* HSPICE Data File for Plotting Id-Vg and Id-Vd Curves in WaveView
.option post=2 ingold=2 numdgt=10

* Independent time source for simulation
VTIME time 0 PWL(0 0 1 1)

* Data table for Id-Vg at Vd = 0.01V
.param vg_data_vd0.01=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.01=[ \
+ 8.817320000000e-11, + 1.286390000000e-10, + 1.876680000000e-10, + 2.737690000000e-10, + 3.993390000000e-10,  \
+ 5.824360000000e-10, + 8.493340000000e-10, + 1.238200000000e-09, + 1.804500000000e-09, + 2.628400000000e-09,  \
+ 3.825400000000e-09, + 5.561200000000e-09, + 8.071600000000e-09, + 1.168790000000e-08, + 1.686830000000e-08,  \
+ 2.423110000000e-08, + 3.458240000000e-08, + 4.892220000000e-08, + 6.840530000000e-08, + 9.423290000000e-08,  \
+ 1.274660000000e-07, + 1.687960000000e-07, + 2.183400000000e-07, + 2.755740000000e-07, + 3.394150000000e-07,  \
+ 4.084390000000e-07, + 4.811210000000e-07, + 5.560310000000e-07, + 6.319470000000e-07, + 7.078840000000e-07,  \
+ 7.830880000000e-07, + 8.570000000000e-07, + 9.292130000000e-07, + 9.994420000000e-07, + 1.067500000000e-06,  \
+ 1.133200000000e-06, + 1.196600000000e-06, + 1.257500000000e-06, + 1.316000000000e-06, + 1.372100000000e-06,  \
+ 1.425800000000e-06, + 1.477200000000e-06, + 1.526300000000e-06, + 1.573200000000e-06, + 1.618000000000e-06,  \
+ 1.660700000000e-06, + 1.701500000000e-06, + 1.740400000000e-06, + 1.777500000000e-06, + 1.812900000000e-06,  \
+ 1.846600000000e-06, + 1.878800000000e-06, + 1.909500000000e-06, + 1.938900000000e-06, + 1.966800000000e-06,  \
+ 1.993600000000e-06, + 2.019100000000e-06, + 2.043500000000e-06, + 2.066800000000e-06, + 2.089000000000e-06,  \
+ 2.110400000000e-06, + 2.130700000000e-06, + 2.150300000000e-06, + 2.168900000000e-06, + 2.186800000000e-06,  \
+ 2.204000000000e-06, + 2.220400000000e-06, + 2.236200000000e-06, + 2.251400000000e-06, + 2.265900000000e-06,  \
+ 2.279900000000e-06, + 2.293300000000e-06, + 2.306100000000e-06, + 2.318500000000e-06, + 2.330500000000e-06,  \
+ 2.341900000000e-06, + 2.353000000000e-06, + 2.363600000000e-06, + 2.373800000000e-06, + 2.383700000000e-06 ]

.param id_pred_data_vd0.01=[ \
+ 8.691662500837e-11, + 1.277592787119e-10, + 1.880239075547e-10, + 2.764217832407e-10, + 4.053875102272e-10,  \
+ 5.927359936209e-10, + 8.640822102279e-10, + 1.256348838297e-09, + 1.822785691274e-09, + 2.640145453370e-09,  \
+ 3.818819322987e-09, + 5.517154022527e-09, + 7.961099299791e-09, + 1.146998670265e-08, + 1.648744500926e-08,  \
+ 2.361348151680e-08, + 3.362896677572e-08, + 4.749799700221e-08, + 6.633278644586e-08, + 9.130706530414e-08,  \
+ 1.235211311723e-07, + 1.638347202970e-07, + 2.127103289240e-07, + 2.701012999751e-07, + 3.354234286235e-07,  \
+ 4.076106051798e-07, + 4.852415804635e-07, + 5.667030200129e-07, + 6.503488111775e-07, + 7.346443453571e-07,  \
+ 8.182539022528e-07, + 9.000972931972e-07, + 9.793627395993e-07, + 1.055493412423e-06, + 1.128153744503e-06,  \
+ 1.197192468680e-06, + 1.262591831619e-06, + 1.324447366642e-06, + 1.382917980663e-06, + 1.438197796233e-06,  \
+ 1.490507129347e-06, + 1.540072262287e-06, + 1.587107253727e-06, + 1.631817576708e-06, + 1.674392406130e-06,  \
+ 1.714990648907e-06, + 1.753766118782e-06, + 1.790846145013e-06, + 1.826332882047e-06, + 1.860323245637e-06,  \
+ 1.892898144433e-06, + 1.924123062054e-06, + 1.954048930202e-06, + 1.982726535061e-06, + 2.010194730246e-06,  \
+ 2.036487130681e-06, + 2.061634586425e-06, + 2.085659943987e-06, + 2.108589542331e-06, + 2.130443899659e-06,  \
+ 2.151242224500e-06, + 2.171011292376e-06, + 2.189765073126e-06, + 2.207524812547e-06, + 2.224314666819e-06,  \
+ 2.240150934085e-06, + 2.255063009216e-06, + 2.269070246257e-06, + 2.282193454448e-06, + 2.294464648003e-06,  \
+ 2.305899979547e-06, + 2.316530444659e-06, + 2.326384565094e-06, + 2.335485332878e-06, + 2.343859378016e-06,  \
+ 2.351536677452e-06, + 2.358541823924e-06, + 2.364902320551e-06, + 2.370651345700e-06, + 2.375804906478e-06 ]

* Data table for Id-Vg at Vd = 0.02V
.param vg_data_vd0.02=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.02=[ \
+ 1.486460000000e-10, + 2.168620000000e-10, + 3.163730000000e-10, + 4.615240000000e-10, + 6.732230000000e-10,  \
+ 9.819230000000e-10, + 1.432000000000e-09, + 2.087800000000e-09, + 3.043000000000e-09, + 4.433200000000e-09,  \
+ 6.454000000000e-09, + 9.386900000000e-09, + 1.363300000000e-08, + 1.975940000000e-08, + 2.855550000000e-08,  \
+ 4.109760000000e-08, + 5.881010000000e-08, + 8.349890000000e-08, + 1.173190000000e-07, + 1.626270000000e-07,  \
+ 2.216860000000e-07, + 2.962440000000e-07, + 3.871040000000e-07, + 4.938470000000e-07, + 6.148470000000e-07,  \
+ 7.475790000000e-07, + 8.890820000000e-07, + 1.036400000000e-06, + 1.186900000000e-06, + 1.338300000000e-06,  \
+ 1.489100000000e-06, + 1.637700000000e-06, + 1.783400000000e-06, + 1.925400000000e-06, + 2.063200000000e-06,  \
+ 2.196600000000e-06, + 2.325300000000e-06, + 2.449200000000e-06, + 2.568300000000e-06, + 2.682600000000e-06,  \
+ 2.792100000000e-06, + 2.896900000000e-06, + 2.997200000000e-06, + 3.093000000000e-06, + 3.184600000000e-06,  \
+ 3.272000000000e-06, + 3.355400000000e-06, + 3.435000000000e-06, + 3.510900000000e-06, + 3.583400000000e-06,  \
+ 3.652500000000e-06, + 3.718400000000e-06, + 3.781300000000e-06, + 3.841400000000e-06, + 3.898700000000e-06,  \
+ 3.953400000000e-06, + 4.005700000000e-06, + 4.055600000000e-06, + 4.103400000000e-06, + 4.149000000000e-06,  \
+ 4.192600000000e-06, + 4.234400000000e-06, + 4.274300000000e-06, + 4.312600000000e-06, + 4.349200000000e-06,  \
+ 4.384300000000e-06, + 4.418000000000e-06, + 4.450300000000e-06, + 4.481200000000e-06, + 4.511000000000e-06,  \
+ 4.539500000000e-06, + 4.566900000000e-06, + 4.593300000000e-06, + 4.618600000000e-06, + 4.642900000000e-06,  \
+ 4.666400000000e-06, + 4.688900000000e-06, + 4.710600000000e-06, + 4.731500000000e-06, + 4.751600000000e-06 ]

.param id_pred_data_vd0.02=[ \
+ 1.456778697673e-10, + 2.137981525152e-10, + 3.144101157204e-10, + 4.621736593435e-10, + 6.780781092175e-10,  \
+ 9.922707278065e-10, + 1.448235451562e-09, + 2.108810548407e-09, + 3.064841394007e-09, + 4.447545052244e-09,  \
+ 6.446107931879e-09, + 9.332759987046e-09, + 1.349756416857e-08, + 1.949491434061e-08, + 2.810066689563e-08,  \
+ 4.037383405375e-08, + 5.770816642325e-08, + 8.184872058337e-08, + 1.148444607679e-07, + 1.589088060427e-07,  \
+ 2.161866723327e-07, + 2.884577588702e-07, + 3.768338865484e-07, + 4.815354259335e-07, + 6.017924533808e-07,  \
+ 7.359194569290e-07, + 8.815071487334e-07, + 1.035695968312e-06, + 1.195480508613e-06, + 1.357968139928e-06,  \
+ 1.520556397736e-06, + 1.681071589701e-06, + 1.837807503762e-06, + 1.989515876630e-06, + 2.135361282853e-06,  \
+ 2.274858561577e-06, + 2.407824067632e-06, + 2.534262021072e-06, + 2.654354320839e-06, + 2.768358681351e-06,  \
+ 2.876606886275e-06, + 2.979459532071e-06, + 3.077284782194e-06, + 3.170417621732e-06, + 3.259199729655e-06,  \
+ 3.343930875417e-06, + 3.424868918955e-06, + 3.502264444251e-06, + 3.576319722924e-06, + 3.647225094028e-06,  \
+ 3.715129569173e-06, + 3.780175466090e-06, + 3.842466685455e-06, + 3.902113239747e-06, + 3.959187888540e-06,  \
+ 4.013780853711e-06, + 4.065953544341e-06, + 4.115761548746e-06, + 4.163260164205e-06, + 4.208500904497e-06,  \
+ 4.251544014551e-06, + 4.292435187381e-06, + 4.331203526817e-06, + 4.367905203253e-06, + 4.402603954077e-06,  \
+ 4.435340233613e-06, + 4.466147220228e-06, + 4.495097091421e-06, + 4.522241652012e-06, + 4.547615535557e-06,  \
+ 4.571282770485e-06, + 4.593307676259e-06, + 4.613730998244e-06, + 4.632619093172e-06, + 4.650023474824e-06,  \
+ 4.666011082008e-06, + 4.680624988396e-06, + 4.693928058259e-06, + 4.705985193141e-06, + 4.716831608675e-06 ]

* Data table for Id-Vg at Vd = 0.03V
.param vg_data_vd0.03=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.03=[ \
+ 1.899920000000e-10, + 2.771750000000e-10, + 4.043540000000e-10, + 5.898610000000e-10, + 8.604170000000e-10,  \
+ 1.255000000000e-09, + 1.830200000000e-09, + 2.668500000000e-09, + 3.889600000000e-09, + 5.667200000000e-09,  \
+ 8.252200000000e-09, + 1.200550000000e-08, + 1.744360000000e-08, + 2.529830000000e-08, + 3.659350000000e-08,  \
+ 5.273540000000e-08, + 7.560430000000e-08, + 1.076220000000e-07, + 1.517480000000e-07, + 2.113360000000e-07,  \
+ 2.898030000000e-07, + 3.900970000000e-07, + 5.140750000000e-07, + 6.619870000000e-07, + 8.322910000000e-07,  \
+ 1.021900000000e-06, + 1.226700000000e-06, + 1.442300000000e-06, + 1.664600000000e-06, + 1.890000000000e-06,  \
+ 2.115400000000e-06, + 2.338800000000e-06, + 2.558400000000e-06, + 2.773000000000e-06, + 2.981800000000e-06,  \
+ 3.184200000000e-06, + 3.379800000000e-06, + 3.568400000000e-06, + 3.749900000000e-06, + 3.924200000000e-06,  \
+ 4.091400000000e-06, + 4.251600000000e-06, + 4.404900000000e-06, + 4.551600000000e-06, + 4.691700000000e-06,  \
+ 4.825600000000e-06, + 4.953500000000e-06, + 5.075600000000e-06, + 5.192100000000e-06, + 5.303300000000e-06,  \
+ 5.409400000000e-06, + 5.510600000000e-06, + 5.607300000000e-06, + 5.699500000000e-06, + 5.787600000000e-06,  \
+ 5.871700000000e-06, + 5.952000000000e-06, + 6.028800000000e-06, + 6.102100000000e-06, + 6.172200000000e-06,  \
+ 6.239300000000e-06, + 6.303500000000e-06, + 6.364900000000e-06, + 6.423700000000e-06, + 6.480000000000e-06,  \
+ 6.533900000000e-06, + 6.585600000000e-06, + 6.635200000000e-06, + 6.682800000000e-06, + 6.728400000000e-06,  \
+ 6.772300000000e-06, + 6.814400000000e-06, + 6.854800000000e-06, + 6.893700000000e-06, + 6.931000000000e-06,  \
+ 6.967000000000e-06, + 7.001500000000e-06, + 7.034800000000e-06, + 7.066900000000e-06, + 7.097700000000e-06 ]

.param id_pred_data_vd0.03=[ \
+ 1.861711851348e-10, + 2.727115866463e-10, + 4.005906539817e-10, + 5.885365261804e-10, + 8.634202686153e-10,  \
+ 1.263943296692e-09, + 1.846051844723e-09, + 2.690773897029e-09, + 3.915456119330e-09, + 5.689836655165e-09,  \
+ 8.259114565590e-09, + 1.197685151055e-08, + 1.735140926939e-08, + 2.510861577321e-08, + 3.627082378443e-08,  \
+ 5.224448159424e-08, + 7.489924200854e-08, + 1.066047593667e-07, + 1.501863380327e-07, + 2.087576285703e-07,  \
+ 2.854238300642e-07, + 3.828816807072e-07, + 5.029957719671e-07, + 6.464607758971e-07, + 8.126270950015e-07,  \
+ 9.995388973039e-07, + 1.204168656841e-06, + 1.422750356141e-06, + 1.651201637287e-06, + 1.885468955152e-06,  \
+ 2.121807192452e-06, + 2.356989207328e-06, + 2.588389324956e-06, + 2.813984756358e-06, + 3.032336171600e-06,  \
+ 3.242508028052e-06, + 3.443980385782e-06, + 3.636576220742e-06, + 3.820327401627e-06, + 3.995483421022e-06,  \
+ 4.162367113167e-06, + 4.321387968957e-06, + 4.472975560930e-06, + 4.617573868018e-06, + 4.755594563903e-06,  \
+ 4.887438408332e-06, + 5.013476475142e-06, + 5.134036618983e-06, + 5.249405221548e-06, + 5.359851638786e-06,  \
+ 5.465596768772e-06, + 5.566840991378e-06, + 5.663767224178e-06, + 5.756525642937e-06, + 5.845231935382e-06,  \
+ 5.930037586950e-06, + 6.011049990775e-06, + 6.088336376706e-06, + 6.162013305584e-06, + 6.232170271687e-06,  \
+ 6.298883672571e-06, + 6.362226413330e-06, + 6.422291044146e-06, + 6.479158764705e-06, + 6.532890693052e-06,  \
+ 6.583595095435e-06, + 6.631333963014e-06, + 6.676190241706e-06, + 6.718261283822e-06, + 6.757625669707e-06,  \
+ 6.794355867896e-06, + 6.828569748905e-06, + 6.860331923235e-06, + 6.889737996971e-06, + 6.916875281604e-06,  \
+ 6.941835017642e-06, + 6.964712374611e-06, + 6.985573272686e-06, + 7.004532089923e-06, + 7.021653873380e-06 ]

* Data table for Id-Vg at Vd = 0.04V
.param vg_data_vd0.04=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.04=[ \
+ 2.183440000000e-10, + 3.185250000000e-10, + 4.646600000000e-10, + 6.778100000000e-10, + 9.886780000000e-10,  \
+ 1.442000000000e-09, + 2.102900000000e-09, + 3.066100000000e-09, + 4.469400000000e-09, + 6.512300000000e-09,  \
+ 9.483700000000e-09, + 1.379950000000e-08, + 2.005540000000e-08, + 2.909780000000e-08, + 4.211440000000e-08,  \
+ 6.074440000000e-08, + 8.719530000000e-08, + 1.243410000000e-07, + 1.757520000000e-07, + 2.455780000000e-07,  \
+ 3.382250000000e-07, + 4.577830000000e-07, + 6.072940000000e-07, + 7.880430000000e-07, + 9.991350000000e-07,  \
+ 1.237500000000e-06, + 1.498600000000e-06, + 1.776700000000e-06, + 2.066400000000e-06, + 2.362500000000e-06,  \
+ 2.660700000000e-06, + 2.957700000000e-06, + 3.250900000000e-06, + 3.538300000000e-06, + 3.818600000000e-06,  \
+ 4.090900000000e-06, + 4.354500000000e-06, + 4.609100000000e-06, + 4.854400000000e-06, + 5.090300000000e-06,  \
+ 5.316800000000e-06, + 5.534000000000e-06, + 5.742200000000e-06, + 5.941400000000e-06, + 6.132000000000e-06,  \
+ 6.314200000000e-06, + 6.488200000000e-06, + 6.654500000000e-06, + 6.813300000000e-06, + 6.964900000000e-06,  \
+ 7.109600000000e-06, + 7.247800000000e-06, + 7.379700000000e-06, + 7.505700000000e-06, + 7.626000000000e-06,  \
+ 7.740800000000e-06, + 7.850600000000e-06, + 7.955500000000e-06, + 8.055700000000e-06, + 8.151600000000e-06,  \
+ 8.243200000000e-06, + 8.331000000000e-06, + 8.414900000000e-06, + 8.495300000000e-06, + 8.572200000000e-06,  \
+ 8.646000000000e-06, + 8.716700000000e-06, + 8.784500000000e-06, + 8.849500000000e-06, + 8.911800000000e-06,  \
+ 8.971700000000e-06, + 9.029200000000e-06, + 9.084400000000e-06, + 9.137500000000e-06, + 9.188500000000e-06,  \
+ 9.237600000000e-06, + 9.284800000000e-06, + 9.330200000000e-06, + 9.373900000000e-06, + 9.416100000000e-06 ]

.param id_pred_data_vd0.04=[ \
+ 2.147539923669e-10, + 3.139287940712e-10, + 4.604901349126e-10, + 6.759600523765e-10, + 9.912714205029e-10,  \
+ 1.451068811775e-09, + 2.120021065366e-09, + 3.091963662882e-09, + 4.502927026806e-09, + 6.549920499310e-09,  \
+ 9.517726198283e-09, + 1.381769607178e-08, + 2.004281441259e-08, + 2.904286247940e-08, + 4.202117906971e-08,  \
+ 6.064481567591e-08, + 8.714865543880e-08, + 1.243966380571e-07, + 1.758481448633e-07, + 2.453843990224e-07,  \
+ 3.369668775122e-07, + 4.541664384305e-07, + 5.996409527143e-07, + 7.746887422400e-07, + 9.789929754334e-07,  \
+ 1.210605914821e-06, + 1.466180547141e-06, + 1.741349988151e-06, + 2.031215262832e-06, + 2.330768329557e-06,  \
+ 2.635279379319e-06, + 2.940545382444e-06, + 3.243032260798e-06, + 3.539928875398e-06, + 3.829123743344e-06,  \
+ 4.109151195735e-06, + 4.379051970318e-06, + 4.638337413780e-06, + 4.886835231446e-06, + 5.124622839503e-06,  \
+ 5.351967993192e-06, + 5.569222266786e-06, + 5.776832695119e-06, + 5.975256790407e-06, + 6.164967198856e-06,  \
+ 6.346412701532e-06, + 6.520015886053e-06, + 6.686164997518e-06, + 6.845245370641e-06, + 6.997558521107e-06,  \
+ 7.143389084376e-06, + 7.283008890226e-06, + 7.416644948535e-06, + 7.544505642727e-06, + 7.666771416552e-06,  \
+ 7.783600012772e-06, + 7.895150920376e-06, + 8.001574897207e-06, + 8.103001164272e-06, + 8.199548465200e-06,  \
+ 8.291330304928e-06, + 8.378471829928e-06, + 8.461105171591e-06, + 8.539339760318e-06, + 8.613269310445e-06,  \
+ 8.683026535437e-06, + 8.748741820455e-06, + 8.810517028905e-06, + 8.868464501575e-06, + 8.922707638703e-06,  \
+ 8.973396616057e-06, + 9.020622237585e-06, + 9.064507903531e-06, + 9.105193894356e-06, + 9.142809431069e-06,  \
+ 9.177447063848e-06, + 9.209263953380e-06, + 9.238345082849e-06, + 9.264849359170e-06, + 9.288860601373e-06 ]

* Data table for Id-Vg at Vd = 0.05V
.param vg_data_vd0.05=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.05=[ \
+ 2.383360000000e-10, + 3.476720000000e-10, + 5.071520000000e-10, + 7.397580000000e-10, + 1.079000000000e-09,  \
+ 1.573700000000e-09, + 2.294800000000e-09, + 3.345900000000e-09, + 4.877100000000e-09, + 7.106500000000e-09,  \
+ 1.034930000000e-08, + 1.506010000000e-08, + 2.189060000000e-08, + 3.176760000000e-08, + 4.599460000000e-08,  \
+ 6.637600000000e-08, + 9.535320000000e-08, + 1.361270000000e-07, + 1.927150000000e-07, + 2.698700000000e-07,  \
+ 3.727770000000e-07, + 5.064870000000e-07, + 6.751480000000e-07, + 8.811830000000e-07, + 1.124700000000e-06,  \
+ 1.403200000000e-06, + 1.712200000000e-06, + 2.045400000000e-06, + 2.396300000000e-06, + 2.758300000000e-06,  \
+ 3.125800000000e-06, + 3.494000000000e-06, + 3.859200000000e-06, + 4.218600000000e-06, + 4.570300000000e-06,  \
+ 4.912800000000e-06, + 5.245000000000e-06, + 5.566400000000e-06, + 5.876600000000e-06, + 6.175300000000e-06,  \
+ 6.462600000000e-06, + 6.738400000000e-06, + 7.002900000000e-06, + 7.256300000000e-06, + 7.498900000000e-06,  \
+ 7.731000000000e-06, + 7.953000000000e-06, + 8.165200000000e-06, + 8.367900000000e-06, + 8.561500000000e-06,  \
+ 8.746500000000e-06, + 8.923200000000e-06, + 9.092000000000e-06, + 9.253200000000e-06, + 9.407200000000e-06,  \
+ 9.554300000000e-06, + 9.694900000000e-06, + 9.829200000000e-06, + 9.957700000000e-06, + 1.008050000000e-05,  \
+ 1.019800000000e-05, + 1.031050000000e-05, + 1.041810000000e-05, + 1.052110000000e-05, + 1.061980000000e-05,  \
+ 1.071440000000e-05, + 1.080500000000e-05, + 1.089190000000e-05, + 1.097520000000e-05, + 1.105520000000e-05,  \
+ 1.113190000000e-05, + 1.120560000000e-05, + 1.127640000000e-05, + 1.134440000000e-05, + 1.140980000000e-05,  \
+ 1.147260000000e-05, + 1.153300000000e-05, + 1.159120000000e-05, + 1.164710000000e-05, + 1.170100000000e-05 ]

.param id_pred_data_vd0.05=[ \
+ 2.355277750610e-10, + 3.435613127323e-10, + 5.031818961498e-10, + 7.378449407014e-10, + 1.081305445183e-09,  \
+ 1.582378850173e-09, + 2.311887747908e-09, + 3.372719703520e-09, + 4.914190654404e-09, + 7.152573999747e-09,  \
+ 1.040068298153e-08, + 1.511071019422e-08, + 2.193568917619e-08, + 3.181422414400e-08, + 4.608139363427e-08,  \
+ 6.659748237325e-08, + 9.587531621946e-08, + 1.371651592308e-07, + 1.944390760400e-07, + 2.722191993598e-07,  \
+ 3.752195880224e-07, + 5.078163667349e-07, + 6.734534963471e-07, + 8.741022611503e-07, + 1.109917866415e-06,  \
+ 1.379164314130e-06, + 1.678416447248e-06, + 2.002974542847e-06, + 2.347348890908e-06, + 2.705799488467e-06,  \
+ 3.072764229728e-06, + 3.443157766014e-06, + 3.812617069343e-06, + 4.177544178674e-06, + 4.535140033113e-06,  \
+ 4.883340807282e-06, + 5.220705497777e-06, + 5.546330430661e-06, + 5.859757584403e-06, + 6.160829070723e-06,  \
+ 6.449643842643e-06, + 6.726470019203e-06, + 6.991661211941e-06, + 7.245667802636e-06, + 7.488935079891e-06,  \
+ 7.721937436145e-06, + 7.945130346343e-06, + 8.158932178048e-06, + 8.363750384888e-06, + 8.559935668018e-06,  \
+ 8.747848914936e-06, + 8.927780436352e-06, + 9.100011084229e-06, + 9.264804975828e-06, + 9.422370203538e-06,  \
+ 9.572932322044e-06, + 9.716676140670e-06, + 9.853797382675e-06, + 9.984461212298e-06, + 1.010882406263e-05,  \
+ 1.022709620884e-05, + 1.033935404848e-05, + 1.044582822942e-05, + 1.054660824593e-05, + 1.064189273166e-05,  \
+ 1.073182502296e-05, + 1.081657319446e-05, + 1.089627403417e-05, + 1.097108906833e-05, + 1.104117181967e-05,  \
+ 1.110668090405e-05, + 1.116779603763e-05, + 1.122467510868e-05, + 1.127743380493e-05, + 1.132628094638e-05,  \
+ 1.137135914178e-05, + 1.141282846220e-05, + 1.145082278526e-05, + 1.148552546510e-05, + 1.151707037934e-05 ]

* Data table for Id-Vg at Vd = 0.06V
.param vg_data_vd0.06=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.06=[ \
+ 2.531020000000e-10, + 3.691890000000e-10, + 5.385060000000e-10, + 7.854450000000e-10, + 1.145600000000e-09,  \
+ 1.670600000000e-09, + 2.436100000000e-09, + 3.551800000000e-09, + 5.177000000000e-09, + 7.543300000000e-09,  \
+ 1.098530000000e-08, + 1.598600000000e-08, + 2.323780000000e-08, + 3.372640000000e-08, + 4.884020000000e-08,  \
+ 7.050410000000e-08, + 1.013310000000e-07, + 1.447610000000e-07, + 2.051410000000e-07, + 2.876720000000e-07,  \
+ 3.981260000000e-07, + 5.423090000000e-07, + 7.252770000000e-07, + 9.504910000000e-07, + 1.219100000000e-06,  \
+ 1.529600000000e-06, + 1.877800000000e-06, + 2.257800000000e-06, + 2.662200000000e-06, + 3.083600000000e-06,  \
+ 3.514900000000e-06, + 3.950300000000e-06, + 4.384600000000e-06, + 4.814100000000e-06, + 5.235900000000e-06,  \
+ 5.647900000000e-06, + 6.048700000000e-06, + 6.437300000000e-06, + 6.813000000000e-06, + 7.175400000000e-06,  \
+ 7.524400000000e-06, + 7.859900000000e-06, + 8.182100000000e-06, + 8.491100000000e-06, + 8.787300000000e-06,  \
+ 9.070900000000e-06, + 9.342300000000e-06, + 9.602000000000e-06, + 9.850200000000e-06, + 1.008760000000e-05,  \
+ 1.031440000000e-05, + 1.053120000000e-05, + 1.073830000000e-05, + 1.093630000000e-05, + 1.112540000000e-05,  \
+ 1.130630000000e-05, + 1.147910000000e-05, + 1.164430000000e-05, + 1.180230000000e-05, + 1.195340000000e-05,  \
+ 1.209800000000e-05, + 1.223640000000e-05, + 1.236890000000e-05, + 1.249570000000e-05, + 1.261720000000e-05,  \
+ 1.273360000000e-05, + 1.284510000000e-05, + 1.295210000000e-05, + 1.305470000000e-05, + 1.315310000000e-05,  \
+ 1.324760000000e-05, + 1.333830000000e-05, + 1.342540000000e-05, + 1.350900000000e-05, + 1.358940000000e-05,  \
+ 1.366670000000e-05, + 1.374110000000e-05, + 1.381250000000e-05, + 1.388130000000e-05, + 1.394760000000e-05 ]

.param id_pred_data_vd0.06=[ \
+ 2.511506735914e-10, + 3.655796465551e-10, + 5.345861353589e-10, + 7.829743253751e-10, + 1.146501560356e-09,  \
+ 1.676932299688e-09, + 2.449504279411e-09, + 3.573605624752e-09, + 5.208061821804e-09, + 7.582889622881e-09,  \
+ 1.103074623643e-08, + 1.603267492101e-08, + 2.328397613383e-08, + 3.378641622476e-08, + 4.896995619674e-08,  \
+ 7.083703394528e-08, + 1.021099569698e-07, + 1.463373337174e-07, + 2.079014166156e-07, + 2.918547852460e-07,  \
+ 4.035554866277e-07, + 5.481073276314e-07, + 7.297013689822e-07, + 9.510032032267e-07, + 1.212725073856e-06,  \
+ 1.513491224614e-06, + 1.849984037108e-06, + 2.217367655248e-06, + 2.609791554278e-06, + 3.020970834768e-06,  \
+ 3.444665344432e-06, + 3.875065594912e-06, + 4.307022609282e-06, + 4.736216214951e-06, + 5.159159190953e-06,  \
+ 5.573164526140e-06, + 5.976271204418e-06, + 6.367145979311e-06, + 6.744912680006e-06, + 7.109163561836e-06,  \
+ 7.459767221007e-06, + 7.796786958352e-06, + 8.120491693262e-06, + 8.431213209406e-06, + 8.729373221286e-06,  \
+ 9.015401301440e-06, + 9.289737499785e-06, + 9.552805277053e-06, + 9.805042936932e-06, + 1.004681456834e-05,  \
+ 1.027851743856e-05, + 1.050046237651e-05, + 1.071297941962e-05, + 1.091634796467e-05, + 1.111084478907e-05,  \
+ 1.129670214141e-05, + 1.147417235188e-05, + 1.164347719168e-05, + 1.180481660413e-05, + 1.195842021843e-05,  \
+ 1.210446003824e-05, + 1.224316132721e-05, + 1.237466902239e-05, + 1.249925378943e-05, + 1.261705270736e-05,  \
+ 1.272827532375e-05, + 1.283310935833e-05, + 1.293176261242e-05, + 1.302444026805e-05, + 1.311130385147e-05,  \
+ 1.319259259617e-05, + 1.326848723693e-05, + 1.333916938165e-05, + 1.340487040579e-05, + 1.346574397758e-05,  \
+ 1.352204504656e-05, + 1.357392029604e-05, + 1.362157665426e-05, + 1.366520446027e-05, + 1.370497047901e-05 ]

* Data table for Id-Vg at Vd = 0.07V
.param vg_data_vd0.07=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.07=[ \
+ 2.644260000000e-10, + 3.856790000000e-10, + 5.625190000000e-10, + 8.204120000000e-10, + 1.196500000000e-09,  \
+ 1.744800000000e-09, + 2.544100000000e-09, + 3.708900000000e-09, + 5.405800000000e-09, + 7.876200000000e-09,  \
+ 1.146990000000e-08, + 1.669080000000e-08, + 2.426260000000e-08, + 3.521550000000e-08, + 5.100170000000e-08,  \
+ 7.363770000000e-08, + 1.058650000000e-07, + 1.513050000000e-07, + 2.145540000000e-07, + 3.011490000000e-07,  \
+ 4.173120000000e-07, + 5.694210000000e-07, + 7.632530000000e-07, + 1.003100000000e-06, + 1.291100000000e-06,  \
+ 1.626600000000e-06, + 2.006400000000e-06, + 2.424700000000e-06, + 2.874400000000e-06, + 3.347500000000e-06,  \
+ 3.836000000000e-06, + 4.332900000000e-06, + 4.831800000000e-06, + 5.327900000000e-06, + 5.817400000000e-06,  \
+ 6.297300000000e-06, + 6.765600000000e-06, + 7.220800000000e-06, + 7.661900000000e-06, + 8.088300000000e-06,  \
+ 8.499600000000e-06, + 8.895700000000e-06, + 9.276500000000e-06, + 9.642300000000e-06, + 9.993300000000e-06,  \
+ 1.032970000000e-05, + 1.065200000000e-05, + 1.096060000000e-05, + 1.125590000000e-05, + 1.153840000000e-05,  \
+ 1.180860000000e-05, + 1.206700000000e-05, + 1.231410000000e-05, + 1.255020000000e-05, + 1.277610000000e-05,  \
+ 1.299200000000e-05, + 1.319850000000e-05, + 1.339590000000e-05, + 1.358480000000e-05, + 1.376550000000e-05,  \
+ 1.393840000000e-05, + 1.410390000000e-05, + 1.426240000000e-05, + 1.441420000000e-05, + 1.455950000000e-05,  \
+ 1.469880000000e-05, + 1.483240000000e-05, + 1.496040000000e-05, + 1.508310000000e-05, + 1.520090000000e-05,  \
+ 1.531400000000e-05, + 1.542250000000e-05, + 1.552670000000e-05, + 1.562680000000e-05, + 1.572300000000e-05,  \
+ 1.581540000000e-05, + 1.590430000000e-05, + 1.598980000000e-05, + 1.607200000000e-05, + 1.615110000000e-05 ]

.param id_pred_data_vd0.07=[ \
+ 2.633494533555e-10, + 3.825738437158e-10, + 5.585687734566e-10, + 8.171192877882e-10, + 1.195418430910e-09,  \
+ 1.747377211814e-09, + 2.551454514332e-09, + 3.721830488246e-09, + 5.424245301811e-09, + 7.898721321453e-09,  \
+ 1.149206738660e-08, + 1.670562255640e-08, + 2.426447622383e-08, + 3.521495955283e-08, + 5.105474315314e-08,  \
+ 7.388982112388e-08, + 1.065985827609e-07, + 1.529590781502e-07, + 2.176764655815e-07, + 3.062376254093e-07,  \
+ 4.245464970154e-07, + 5.783459801023e-07, + 7.725201703579e-07, + 1.010416999634e-06, + 1.293344266742e-06,  \
+ 1.620377115614e-06, + 1.988452131627e-06, + 2.392755377514e-06, + 2.827268253895e-06, + 3.285329657956e-06,  \
+ 3.760185027204e-06, + 4.245406271366e-06, + 4.735198890558e-06, + 5.224554261076e-06, + 5.709332908737e-06,  \
+ 6.186244136188e-06, + 6.652783122263e-06, + 7.107121418812e-06, + 7.548015273642e-06, + 7.974672698765e-06,  \
+ 8.386695408262e-06, + 8.783935190877e-06, + 9.166457748506e-06, + 9.534508571960e-06, + 9.888352506096e-06,  \
+ 1.022838987410e-05, + 1.055498636561e-05, + 1.086859221687e-05, + 1.116956089390e-05, + 1.145832429756e-05,  \
+ 1.173523080070e-05, + 1.200064201839e-05, + 1.225489817443e-05, + 1.249832013855e-05, + 1.273117377423e-05,  \
+ 1.295377893257e-05, + 1.316638212302e-05, + 1.336925939540e-05, + 1.356264605420e-05, + 1.374678962748e-05,  \
+ 1.392190402839e-05, + 1.408826836268e-05, + 1.424610061804e-05, + 1.439560655854e-05, + 1.453708566260e-05,  \
+ 1.467068970669e-05, + 1.479671409470e-05, + 1.491536866524e-05, + 1.502690502093e-05, + 1.513155235443e-05,  \
+ 1.522954902612e-05, + 1.532113543362e-05, + 1.540652854601e-05, + 1.548602987896e-05, + 1.555976676173e-05,  \
+ 1.562808654853e-05, + 1.569113897858e-05, + 1.574921741849e-05, + 1.580249198014e-05, + 1.585118370713e-05 ]

* Data table for Id-Vg at Vd = 0.08V
.param vg_data_vd0.08=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.08=[ \
+ 2.733620000000e-10, + 3.986810000000e-10, + 5.814360000000e-10, + 8.479340000000e-10, + 1.236500000000e-09,  \
+ 1.803000000000e-09, + 2.628800000000e-09, + 3.832200000000e-09, + 5.585100000000e-09, + 8.137000000000e-09,  \
+ 1.184890000000e-08, + 1.724170000000e-08, + 2.506280000000e-08, + 3.637710000000e-08, + 5.268640000000e-08,  \
+ 7.607750000000e-08, + 1.093920000000e-07, + 1.563890000000e-07, + 2.218590000000e-07, + 3.115980000000e-07,  \
+ 4.321700000000e-07, + 5.904030000000e-07, + 7.926320000000e-07, + 1.043800000000e-06, + 1.346900000000e-06,  \
+ 1.702100000000e-06, + 2.106900000000e-06, + 2.556400000000e-06, + 3.043600000000e-06, + 3.560600000000e-06,  \
+ 4.099000000000e-06, + 4.650600000000e-06, + 5.208500000000e-06, + 5.766500000000e-06, + 6.319800000000e-06,  \
+ 6.864700000000e-06, + 7.398400000000e-06, + 7.918700000000e-06, + 8.424300000000e-06, + 8.914200000000e-06,  \
+ 9.387800000000e-06, + 9.844600000000e-06, + 1.028470000000e-05, + 1.070800000000e-05, + 1.111460000000e-05,  \
+ 1.150500000000e-05, + 1.187930000000e-05, + 1.223810000000e-05, + 1.258180000000e-05, + 1.291080000000e-05,  \
+ 1.322580000000e-05, + 1.352720000000e-05, + 1.381560000000e-05, + 1.409140000000e-05, + 1.435530000000e-05,  \
+ 1.460770000000e-05, + 1.484920000000e-05, + 1.508020000000e-05, + 1.530130000000e-05, + 1.551280000000e-05,  \
+ 1.571530000000e-05, + 1.590920000000e-05, + 1.609480000000e-05, + 1.627260000000e-05, + 1.644300000000e-05,  \
+ 1.660620000000e-05, + 1.676270000000e-05, + 1.691270000000e-05, + 1.705660000000e-05, + 1.719470000000e-05,  \
+ 1.732710000000e-05, + 1.745430000000e-05, + 1.757640000000e-05, + 1.769370000000e-05, + 1.780640000000e-05,  \
+ 1.791470000000e-05, + 1.801870000000e-05, + 1.811880000000e-05, + 1.821510000000e-05, + 1.830770000000e-05 ]

.param id_pred_data_vd0.08=[ \
+ 2.732483928014e-10, + 3.962265537893e-10, + 5.776620071174e-10, + 8.440661503073e-10, + 1.233691904190e-09,  \
+ 1.802077918001e-09, + 2.630122253322e-09, + 3.835617974346e-09, + 5.589569127551e-09, + 8.139339229274e-09,  \
+ 1.184209281746e-08, + 1.721363787510e-08, + 2.499994707250e-08, + 3.627864316513e-08, + 5.259542376734e-08,  \
+ 7.613099114678e-08, + 1.098793109122e-07, + 1.577928196639e-07, + 2.248303098895e-07, + 3.168278999510e-07,  \
+ 4.401463957038e-07, + 6.010840661475e-07, + 8.051475015236e-07, + 1.056331748259e-06, + 1.356550783385e-06,  \
+ 1.705380127532e-06, + 2.100105484715e-06, + 2.536080137361e-06, + 3.007243794855e-06, + 3.506719367579e-06,  \
+ 4.027392715216e-06, + 4.562345857266e-06, + 5.105215823278e-06, + 5.650414386764e-06, + 6.193214212544e-06,  \
+ 6.729720043950e-06, + 7.256902172230e-06, + 7.772432873026e-06, + 8.274642750621e-06, + 8.762364741415e-06,  \
+ 9.234870085493e-06, + 9.691776940599e-06, + 1.013291068375e-05, + 1.055830740370e-05, + 1.096818596125e-05,  \
+ 1.136274659075e-05, + 1.174232689664e-05, + 1.210729475133e-05, + 1.245797728188e-05, + 1.279478077777e-05,  \
+ 1.311803935096e-05, + 1.342811272480e-05, + 1.372536877170e-05, + 1.401007291861e-05, + 1.428260933608e-05,  \
+ 1.454325392842e-05, + 1.479228143580e-05, + 1.503001200035e-05, + 1.525667263195e-05, + 1.547260791995e-05,  \
+ 1.567804836668e-05, + 1.587329781614e-05, + 1.605861471035e-05, + 1.623423187993e-05, + 1.640047412366e-05,  \
+ 1.655759755522e-05, + 1.670588389970e-05, + 1.684556598775e-05, + 1.697700703517e-05, + 1.710038864985e-05,  \
+ 1.721607754007e-05, + 1.732428558171e-05, + 1.742531196214e-05, + 1.751944073476e-05, + 1.760693965480e-05,  \
+ 1.768811140209e-05, + 1.776316668838e-05, + 1.783241750672e-05, + 1.789610134438e-05, + 1.795449759811e-05 ]

* Data table for Id-Vg at Vd = 0.09V
.param vg_data_vd0.09=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.09=[ \
+ 2.806440000000e-10, + 4.092660000000e-10, + 5.968220000000e-10, + 8.702980000000e-10, + 1.269000000000e-09,  \
+ 1.850300000000e-09, + 2.697500000000e-09, + 3.931900000000e-09, + 5.730000000000e-09, + 8.347500000000e-09,  \
+ 1.215470000000e-08, + 1.768560000000e-08, + 2.570680000000e-08, + 3.731070000000e-08, + 5.403840000000e-08,  \
+ 7.803240000000e-08, + 1.122130000000e-07, + 1.604480000000e-07, + 2.276780000000e-07, + 3.199010000000e-07,  \
+ 4.439490000000e-07, + 6.069940000000e-07, + 8.158120000000e-07, + 1.075900000000e-06, + 1.390900000000e-06,  \
+ 1.761600000000e-06, + 2.186400000000e-06, + 2.661000000000e-06, + 3.179000000000e-06, + 3.732700000000e-06,  \
+ 4.313500000000e-06, + 4.913100000000e-06, + 5.523500000000e-06, + 6.137900000000e-06, + 6.750400000000e-06,  \
+ 7.356300000000e-06, + 7.952200000000e-06, + 8.535200000000e-06, + 9.103500000000e-06, + 9.655600000000e-06,  \
+ 1.019060000000e-05, + 1.070780000000e-05, + 1.120700000000e-05, + 1.168790000000e-05, + 1.215080000000e-05,  \
+ 1.259560000000e-05, + 1.302290000000e-05, + 1.343280000000e-05, + 1.382590000000e-05, + 1.420270000000e-05,  \
+ 1.456360000000e-05, + 1.490930000000e-05, + 1.524030000000e-05, + 1.555710000000e-05, + 1.586030000000e-05,  \
+ 1.615050000000e-05, + 1.642830000000e-05, + 1.669420000000e-05, + 1.694870000000e-05, + 1.719230000000e-05,  \
+ 1.742560000000e-05, + 1.764890000000e-05, + 1.786290000000e-05, + 1.806780000000e-05, + 1.826420000000e-05,  \
+ 1.845240000000e-05, + 1.863290000000e-05, + 1.880590000000e-05, + 1.897180000000e-05, + 1.913100000000e-05,  \
+ 1.928380000000e-05, + 1.943040000000e-05, + 1.957120000000e-05, + 1.970640000000e-05, + 1.983630000000e-05,  \
+ 1.996110000000e-05, + 2.008100000000e-05, + 2.019630000000e-05, + 2.030720000000e-05, + 2.041390000000e-05 ]

.param id_pred_data_vd0.09=[ \
+ 2.815800392852e-10, + 4.076364046313e-10, + 5.935148772451e-10, + 8.662843242746e-10, + 1.265036475573e-09,  \
+ 1.846566899388e-09, + 2.693707017443e-09, + 3.927132858905e-09, + 5.721949634108e-09, + 8.331265277661e-09,  \
+ 1.211989740568e-08, + 1.761427739666e-08, + 2.557515159651e-08, + 3.710213064778e-08, + 5.377482011681e-08,  \
+ 7.782760803821e-08, + 1.123392758018e-07, + 1.613942515633e-07, + 2.301471704413e-07, + 3.247158906561e-07,  \
+ 4.518352898231e-07, + 6.182780316522e-07, + 8.301041543746e-07, + 1.091902831831e-06, + 1.406178034813e-06,  \
+ 1.773029871401e-06, + 2.190153481934e-06, + 2.653153278516e-06, + 3.156062557537e-06, + 3.691908787005e-06,  \
+ 4.253350271028e-06, + 4.833094753849e-06, + 5.424353548733e-06, + 6.021007211530e-06, + 6.617785620620e-06,  \
+ 7.210285330075e-06, + 7.794950579409e-06, + 8.368976050406e-06, + 8.930241383496e-06, + 9.477190033067e-06,  \
+ 1.000876181934e-05, + 1.052426261595e-05, + 1.102326481487e-05, + 1.150565381977e-05, + 1.197134843096e-05,  \
+ 1.242053069291e-05, + 1.285341670155e-05, + 1.327022124315e-05, + 1.367123899399e-05, + 1.405684059137e-05,  \
+ 1.442729058908e-05, + 1.478297926951e-05, + 1.512419868959e-05, + 1.545129198348e-05, + 1.576459442731e-05,  \
+ 1.606436664588e-05, + 1.635095963138e-05, + 1.662467591814e-05, + 1.688583244686e-05, + 1.713474353892e-05,  \
+ 1.737165934173e-05, + 1.759692691849e-05, + 1.781084094546e-05, + 1.801371050533e-05, + 1.820584599045e-05,  \
+ 1.838754207711e-05, + 1.855911832536e-05, + 1.872091917903e-05, + 1.887325634016e-05, + 1.901640091091e-05,  \
+ 1.915071305120e-05, + 1.927648481796e-05, + 1.939409208717e-05, + 1.950374833541e-05, + 1.960590670933e-05,  \
+ 1.970074532437e-05, + 1.978864398552e-05, + 1.986990260775e-05, + 1.994479884161e-05, + 2.001362081501e-05 ]

* Data table for Id-Vg at Vd = 0.10V
.param vg_data_vd0.10=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.10=[ \
+ 2.868030000000e-10, + 4.182090000000e-10, + 6.098080000000e-10, + 8.891530000000e-10, + 1.296400000000e-09,  \
+ 1.890000000000e-09, + 2.755200000000e-09, + 4.015700000000e-09, + 5.851500000000e-09, + 8.523800000000e-09,  \
+ 1.241040000000e-08, + 1.805630000000e-08, + 2.624390000000e-08, + 3.808810000000e-08, + 5.516210000000e-08,  \
+ 7.965400000000e-08, + 1.145470000000e-07, + 1.637980000000e-07, + 2.324640000000e-07, + 3.267040000000e-07,  \
+ 4.535590000000e-07, + 6.204690000000e-07, + 8.345510000000e-07, + 1.101800000000e-06, + 1.426100000000e-06,  \
+ 1.809200000000e-06, + 2.249900000000e-06, + 2.744700000000e-06, + 3.287800000000e-06, + 3.871800000000e-06,  \
+ 4.488500000000e-06, + 5.129300000000e-06, + 5.785900000000e-06, + 6.450700000000e-06, + 7.117000000000e-06,  \
+ 7.779500000000e-06, + 8.433700000000e-06, + 9.076200000000e-06, + 9.704600000000e-06, + 1.031680000000e-05,  \
+ 1.091160000000e-05, + 1.148810000000e-05, + 1.204560000000e-05, + 1.258380000000e-05, + 1.310270000000e-05,  \
+ 1.360230000000e-05, + 1.408280000000e-05, + 1.454450000000e-05, + 1.498780000000e-05, + 1.541310000000e-05,  \
+ 1.582100000000e-05, + 1.621200000000e-05, + 1.658660000000e-05, + 1.694560000000e-05, + 1.728930000000e-05,  \
+ 1.761850000000e-05, + 1.793380000000e-05, + 1.823570000000e-05, + 1.852480000000e-05, + 1.880170000000e-05,  \
+ 1.906680000000e-05, + 1.932080000000e-05, + 1.956420000000e-05, + 1.979730000000e-05, + 2.002080000000e-05,  \
+ 2.023500000000e-05, + 2.044030000000e-05, + 2.063720000000e-05, + 2.082610000000e-05, + 2.100730000000e-05,  \
+ 2.118120000000e-05, + 2.134810000000e-05, + 2.150830000000e-05, + 2.166220000000e-05, + 2.180990000000e-05,  \
+ 2.195190000000e-05, + 2.208840000000e-05, + 2.221950000000e-05, + 2.234560000000e-05, + 2.246680000000e-05 ]

.param id_pred_data_vd0.10=[ \
+ 2.888212113916e-10, + 4.175175760679e-10, + 6.071995350965e-10, + 8.853931809938e-10, + 1.291863949149e-09,  \
+ 1.884461120483e-09, + 2.747617777743e-09, + 4.004414932979e-09, + 5.833383909248e-09, + 8.492235537005e-09,  \
+ 1.235191149362e-08, + 1.794673067934e-08, + 2.604829489883e-08, + 3.777169581554e-08, + 5.472063548950e-08,  \
+ 7.916808044683e-08, + 1.142550900113e-07, + 1.641640210437e-07, + 2.342020252399e-07, + 3.307080305603e-07,  \
+ 4.607256414602e-07, + 6.314235179161e-07, + 8.493442692270e-07, + 1.119615080825e-06, + 1.445293219149e-06,  \
+ 1.826999141485e-06, + 2.262871385028e-06, + 2.748838232947e-06, + 3.279096927145e-06, + 3.846712206723e-06,  \
+ 4.444202204468e-06, + 5.064051947556e-06, + 5.699104804080e-06, + 6.342821870930e-06, + 6.989484973019e-06,  \
+ 7.634205394424e-06, + 8.272930426756e-06, + 8.902414265322e-06, + 9.520095773041e-06, + 1.012405264191e-05,  \
+ 1.071283040801e-05, + 1.128541116486e-05, + 1.184113934869e-05, + 1.237961987499e-05, + 1.290061627515e-05,  \
+ 1.340410963167e-05, + 1.389013923472e-05, + 1.435891317669e-05, + 1.481056096964e-05, + 1.524537074147e-05,  \
+ 1.566361024743e-05, + 1.606558362255e-05, + 1.645154115977e-05, + 1.682185393292e-05, + 1.717678242130e-05,  \
+ 1.751671661623e-05, + 1.784185878932e-05, + 1.815264695324e-05, + 1.844930957304e-05, + 1.873221481219e-05,  \
+ 1.900169008877e-05, + 1.925804681377e-05, + 1.950167352334e-05, + 1.973283360712e-05, + 1.995192287723e-05,  \
+ 2.015925274463e-05, + 2.035520155914e-05, + 2.054010401480e-05, + 2.071433409583e-05, + 2.087821194436e-05,  \
+ 2.103213191731e-05, + 2.117643889505e-05, + 2.131151122740e-05, + 2.143770980183e-05, + 2.155532274628e-05,  \
+ 2.166475605918e-05, + 2.176633570343e-05, + 2.186044730479e-05, + 2.194732514909e-05, + 2.202742616646e-05 ]

* Data table for Id-Vg at Vd = 0.11V
.param vg_data_vd0.11=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.11=[ \
+ 2.922060000000e-10, + 4.260460000000e-10, + 6.211740000000e-10, + 9.056390000000e-10, + 1.320300000000e-09,  \
+ 1.924700000000e-09, + 2.805400000000e-09, + 4.088600000000e-09, + 5.957200000000e-09, + 8.676900000000e-09,  \
+ 1.263210000000e-08, + 1.837730000000e-08, + 2.670820000000e-08, + 3.875900000000e-08, + 5.613010000000e-08,  \
+ 8.104760000000e-08, + 1.165480000000e-07, + 1.666590000000e-07, + 2.365380000000e-07, + 3.324680000000e-07,  \
+ 4.616560000000e-07, + 6.317530000000e-07, + 8.501400000000e-07, + 1.123100000000e-06, + 1.455100000000e-06,  \
+ 1.848100000000e-06, + 2.301600000000e-06, + 2.812600000000e-06, + 3.376100000000e-06, + 3.985000000000e-06,  \
+ 4.631600000000e-06, + 5.307400000000e-06, + 6.003900000000e-06, + 6.713100000000e-06, + 7.427800000000e-06,  \
+ 8.141800000000e-06, + 8.850000000000e-06, + 9.548400000000e-06, + 1.023360000000e-05, + 1.090330000000e-05,  \
+ 1.155580000000e-05, + 1.218970000000e-05, + 1.280430000000e-05, + 1.339880000000e-05, + 1.397310000000e-05,  \
+ 1.452710000000e-05, + 1.506070000000e-05, + 1.557430000000e-05, + 1.606810000000e-05, + 1.654250000000e-05,  \
+ 1.699790000000e-05, + 1.743500000000e-05, + 1.785420000000e-05, + 1.825610000000e-05, + 1.864140000000e-05,  \
+ 1.901060000000e-05, + 1.936450000000e-05, + 1.970340000000e-05, + 2.002820000000e-05, + 2.033940000000e-05,  \
+ 2.063750000000e-05, + 2.092320000000e-05, + 2.119690000000e-05, + 2.145930000000e-05, + 2.171080000000e-05,  \
+ 2.195190000000e-05, + 2.218300000000e-05, + 2.240470000000e-05, + 2.261740000000e-05, + 2.282140000000e-05,  \
+ 2.301720000000e-05, + 2.320510000000e-05, + 2.338550000000e-05, + 2.355870000000e-05, + 2.372510000000e-05,  \
+ 2.388490000000e-05, + 2.403840000000e-05, + 2.418600000000e-05, + 2.432780000000e-05, + 2.446420000000e-05 ]

.param id_pred_data_vd0.11=[ \
+ 2.952820987723e-10, + 4.263325914522e-10, + 6.194069834820e-10, + 9.024289759907e-10, + 1.315746560593e-09,  \
+ 1.918109795440e-09, + 2.795372129327e-09, + 4.072723029935e-09, + 5.931702666828e-09, + 8.634034074362e-09,  \
+ 1.255567831038e-08, + 1.823736724305e-08, + 2.645884705998e-08, + 3.834654052071e-08, + 5.552159393574e-08,  \
+ 8.028475690480e-08, + 1.158222596587e-07, + 1.663911734795e-07, + 2.374140058237e-07, + 3.354043860782e-07,  \
+ 4.676530761571e-07, + 6.416612313842e-07, + 8.643805631436e-07, + 1.141416660175e-06, + 1.476336756241e-06,  \
+ 1.870266150945e-06, + 2.321784213564e-06, + 2.827183998306e-06, + 3.380906236998e-06, + 3.976120096922e-06,  \
+ 4.605325448210e-06, + 5.260851685307e-06, + 5.935293520452e-06, + 6.621778302360e-06, + 7.314208924072e-06,  \
+ 8.007257420104e-06, + 8.696480217623e-06, + 9.378142058267e-06, + 1.004934805678e-05, + 1.070771315426e-05,  \
+ 1.135148137109e-05, + 1.197927929752e-05, + 1.259019372810e-05, + 1.318349233770e-05, + 1.375882697175e-05,  \
+ 1.431595112081e-05, + 1.485472152126e-05, + 1.537515738164e-05, + 1.587741397088e-05, + 1.636155851884e-05,  \
+ 1.682783913566e-05, + 1.727650393150e-05, + 1.770773858880e-05, + 1.812189366319e-05, + 1.851922206697e-05,  \
+ 1.890002953587e-05, + 1.926462180563e-05, + 1.961328380276e-05, + 1.994642530917e-05, + 2.026430243859e-05,  \
+ 2.056732977508e-05, + 2.085580345010e-05, + 2.113008042215e-05, + 2.139055446605e-05, + 2.163762255805e-05,  \
+ 2.187160323956e-05, + 2.209291749750e-05, + 2.230191908893e-05, + 2.249903220218e-05, + 2.268468582770e-05,  \
+ 2.285918089910e-05, + 2.302298322320e-05, + 2.317644175491e-05, + 2.332002230105e-05, + 2.345404340304e-05,  \
+ 2.357891804422e-05, + 2.369507681578e-05, + 2.380283825914e-05, + 2.390261055552e-05, + 2.399474426056e-05 ]

* Data table for Id-Vg at Vd = 0.12V
.param vg_data_vd0.12=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.12=[ \
+ 2.970960000000e-10, + 4.331320000000e-10, + 6.314420000000e-10, + 9.205150000000e-10, + 1.341900000000e-09,  \
+ 1.955900000000e-09, + 2.850700000000e-09, + 4.154000000000e-09, + 6.052000000000e-09, + 8.814100000000e-09,  \
+ 1.283060000000e-08, + 1.866420000000e-08, + 2.712270000000e-08, + 3.935690000000e-08, + 5.699100000000e-08,  \
+ 8.228430000000e-08, + 1.183180000000e-07, + 1.691840000000e-07, + 2.401160000000e-07, + 3.375060000000e-07,  \
+ 4.686930000000e-07, + 6.414950000000e-07, + 8.634970000000e-07, + 1.141200000000e-06, + 1.479400000000e-06,  \
+ 1.880600000000e-06, + 2.344500000000e-06, + 2.868800000000e-06, + 3.448800000000e-06, + 4.078200000000e-06,  \
+ 4.749500000000e-06, + 5.454600000000e-06, + 6.185100000000e-06, + 6.932800000000e-06, + 7.690300000000e-06,  \
+ 8.450800000000e-06, + 9.208400000000e-06, + 9.958400000000e-06, + 1.069700000000e-05, + 1.142120000000e-05,  \
+ 1.212880000000e-05, + 1.281800000000e-05, + 1.348770000000e-05, + 1.413710000000e-05, + 1.476560000000e-05,  \
+ 1.537310000000e-05, + 1.595930000000e-05, + 1.652440000000e-05, + 1.706860000000e-05, + 1.759220000000e-05,  \
+ 1.809550000000e-05, + 1.857900000000e-05, + 1.904340000000e-05, + 1.948900000000e-05, + 1.991650000000e-05,  \
+ 2.032660000000e-05, + 2.071980000000e-05, + 2.109680000000e-05, + 2.145810000000e-05, + 2.180460000000e-05,  \
+ 2.213660000000e-05, + 2.245490000000e-05, + 2.276000000000e-05, + 2.305250000000e-05, + 2.333290000000e-05,  \
+ 2.360180000000e-05, + 2.385970000000e-05, + 2.410700000000e-05, + 2.434420000000e-05, + 2.457190000000e-05,  \
+ 2.479030000000e-05, + 2.500000000000e-05, + 2.520120000000e-05, + 2.539450000000e-05, + 2.558000000000e-05,  \
+ 2.575830000000e-05, + 2.592950000000e-05, + 2.609400000000e-05, + 2.625210000000e-05, + 2.640400000000e-05 ]

.param id_pred_data_vd0.12=[ \
+ 3.011657589980e-10, + 4.343790394046e-10, + 6.305873156975e-10, + 9.180662630115e-10, + 1.337685695546e-09,  \
+ 1.949021850578e-09, + 2.839225174966e-09, + 4.135463171906e-09, + 6.022046221688e-09, + 8.764331766997e-09,  \
+ 1.274283675912e-08, + 1.850365833889e-08, + 2.683318143681e-08, + 3.886673766829e-08, + 5.623829679280e-08,  \
+ 8.126902457661e-08, + 1.171790472654e-07, + 1.682807851466e-07, + 2.400854555162e-07, + 3.392421967874e-07,  \
+ 4.732409979624e-07, + 6.498524453491e-07, + 8.763780715526e-07, + 1.158834238595e-06, + 1.501248407294e-06,  \
+ 1.905216195155e-06, + 2.369764188188e-06, + 2.891561016440e-06, + 3.465326080914e-06, + 4.084414104000e-06,  \
+ 4.741357115563e-06, + 5.428439180832e-06, + 6.138083408587e-06, + 6.863198359497e-06, + 7.597338699270e-06,  \
+ 8.334842277691e-06, + 9.070867672563e-06, + 9.801345295273e-06, + 1.052291278029e-05, + 1.123288355302e-05,  \
+ 1.192910625832e-05, + 1.260994904442e-05, + 1.327412581304e-05, + 1.392070669681e-05, + 1.454907964217e-05,  \
+ 1.515874697361e-05, + 1.574943889864e-05, + 1.632103929296e-05, + 1.687349402346e-05, + 1.740682579111e-05,  \
+ 1.792117254809e-05, + 1.841661287472e-05, + 1.889345236123e-05, + 1.935186737683e-05, + 1.979206921533e-05,  \
+ 2.021435124334e-05, + 2.061900158878e-05, + 2.100637299009e-05, + 2.137670817319e-05, + 2.173043321818e-05,  \
+ 2.206783974543e-05, + 2.238929271698e-05, + 2.269524615258e-05, + 2.298599516507e-05, + 2.326196059585e-05,  \
+ 2.352353185415e-05, + 2.377119439188e-05, + 2.400531840976e-05, + 2.422628807835e-05, + 2.443458361086e-05,  \
+ 2.463061886374e-05, + 2.481485134922e-05, + 2.498771063983e-05, + 2.514956169762e-05, + 2.530090219807e-05,  \
+ 2.544218266848e-05, + 2.557371568400e-05, + 2.569604956079e-05, + 2.580946544185e-05, + 2.591446100269e-05 ]

* Data table for Id-Vg at Vd = 0.13V
.param vg_data_vd0.13=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.13=[ \
+ 3.016350000000e-10, + 4.397030000000e-10, + 6.409550000000e-10, + 9.342860000000e-10, + 1.361800000000e-09,  \
+ 1.984800000000e-09, + 2.892400000000e-09, + 4.214400000000e-09, + 6.139300000000e-09, + 8.940300000000e-09,  \
+ 1.301300000000e-08, + 1.892760000000e-08, + 2.750250000000e-08, + 3.990390000000e-08, + 5.777730000000e-08,  \
+ 8.341130000000e-08, + 1.199280000000e-07, + 1.714710000000e-07, + 2.433460000000e-07, + 3.420330000000e-07,  \
+ 4.749800000000e-07, + 6.501380000000e-07, + 8.752560000000e-07, + 1.157100000000e-06, + 1.500500000000e-06,  \
+ 1.908400000000e-06, + 2.381000000000e-06, + 2.916100000000e-06, + 3.509700000000e-06, + 4.155800000000e-06,  \
+ 4.847600000000e-06, + 5.577100000000e-06, + 6.336400000000e-06, + 7.117200000000e-06, + 7.912000000000e-06,  \
+ 8.713600000000e-06, + 9.515700000000e-06, + 1.031310000000e-05, + 1.110120000000e-05, + 1.187650000000e-05,  \
+ 1.263630000000e-05, + 1.337830000000e-05, + 1.410110000000e-05, + 1.480350000000e-05, + 1.548470000000e-05,  \
+ 1.614440000000e-05, + 1.678230000000e-05, + 1.739820000000e-05, + 1.799220000000e-05, + 1.856470000000e-05,  \
+ 1.911570000000e-05, + 1.964590000000e-05, + 2.015550000000e-05, + 2.064520000000e-05, + 2.111550000000e-05,  \
+ 2.156690000000e-05, + 2.200020000000e-05, + 2.241580000000e-05, + 2.281460000000e-05, + 2.319700000000e-05,  \
+ 2.356380000000e-05, + 2.391550000000e-05, + 2.425280000000e-05, + 2.457620000000e-05, + 2.488640000000e-05,  \
+ 2.518390000000e-05, + 2.546920000000e-05, + 2.574300000000e-05, + 2.600560000000e-05, + 2.625760000000e-05,  \
+ 2.649940000000e-05, + 2.673150000000e-05, + 2.695420000000e-05, + 2.716810000000e-05, + 2.737350000000e-05,  \
+ 2.757070000000e-05, + 2.776020000000e-05, + 2.794220000000e-05, + 2.811700000000e-05, + 2.828500000000e-05 ]

.param id_pred_data_vd0.13=[ \
+ 3.066067399971e-10, + 4.418489818470e-10, + 6.410179986815e-10, + 9.327219041566e-10, + 1.358314332123e-09,  \
+ 1.978142236680e-09, + 2.880601872590e-09, + 4.194753842057e-09, + 6.107592867011e-09, + 8.887953057979e-09,  \
+ 1.292070187731e-08, + 1.875687033248e-08, + 2.718873361118e-08, + 3.935887576745e-08, + 5.691141325315e-08,  \
+ 8.218355389999e-08, + 1.184208628047e-07, + 1.699775623365e-07, + 2.424329375117e-07, + 3.425409090596e-07,  \
+ 4.779484288520e-07, + 6.566435104105e-07, + 8.862206095728e-07, + 1.173047648990e-06, + 1.521558533568e-06,  \
+ 1.933775956786e-06, + 2.409151311440e-06, + 2.944735952042e-06, + 3.535564155754e-06, + 4.175199719612e-06,  \
+ 4.856294617639e-06, + 5.571147303272e-06, + 6.312094301393e-06, + 7.071859945427e-06, + 7.843790008337e-06,  \
+ 8.621909873909e-06, + 9.401065472048e-06, + 1.017683767714e-05, + 1.094553001167e-05, + 1.170408824692e-05,  \
+ 1.245005310921e-05, + 1.318145434198e-05, + 1.389674922393e-05, + 1.459472892748e-05, + 1.527450433059e-05,  \
+ 1.593537643203e-05, + 1.657694985624e-05, + 1.719879423035e-05, + 1.780082820915e-05, + 1.838286829297e-05,  \
+ 1.894498069305e-05, + 1.948718811036e-05, + 2.000963810133e-05, + 2.051242146990e-05, + 2.099577468471e-05,  \
+ 2.145996259060e-05, + 2.190518760472e-05, + 2.233179780887e-05, + 2.274006939842e-05, + 2.313031262020e-05,  \
+ 2.350289825699e-05, + 2.385817628237e-05, + 2.419652315439e-05, + 2.451842694427e-05, + 2.482419789885e-05,  \
+ 2.511432598112e-05, + 2.538921980886e-05, + 2.564933151007e-05, + 2.589508862002e-05, + 2.612704920466e-05,  \
+ 2.634552918607e-05, + 2.655112257344e-05, + 2.674423609278e-05, + 2.692529538763e-05, + 2.709489257541e-05,  \
+ 2.725338898017e-05, + 2.740123483818e-05, + 2.753892767942e-05, + 2.766694233287e-05, + 2.778564012260e-05 ]

* Data table for Id-Vg at Vd = 0.14V
.param vg_data_vd0.14=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.14=[ \
+ 3.059300000000e-10, + 4.459170000000e-10, + 6.499420000000e-10, + 9.472830000000e-10, + 1.380600000000e-09,  \
+ 2.011900000000e-09, + 2.931700000000e-09, + 4.271200000000e-09, + 6.221300000000e-09, + 9.058800000000e-09,  \
+ 1.318400000000e-08, + 1.917420000000e-08, + 2.785770000000e-08, + 4.041480000000e-08, + 5.851040000000e-08,  \
+ 8.446020000000e-08, + 1.214220000000e-07, + 1.735890000000e-07, + 2.463260000000e-07, + 3.461910000000e-07,  \
+ 4.807240000000e-07, + 6.579870000000e-07, + 8.858570000000e-07, + 1.171200000000e-06, + 1.519200000000e-06,  \
+ 1.932900000000e-06, + 2.412700000000e-06, + 2.956900000000e-06, + 3.561700000000e-06, + 4.221800000000e-06,  \
+ 4.930400000000e-06, + 5.680400000000e-06, + 6.463700000000e-06, + 7.272700000000e-06, + 8.099600000000e-06,  \
+ 8.937200000000e-06, + 9.779000000000e-06, + 1.061910000000e-05, + 1.145260000000e-05, + 1.227540000000e-05,  \
+ 1.308410000000e-05, + 1.387620000000e-05, + 1.464960000000e-05, + 1.540300000000e-05, + 1.613520000000e-05,  \
+ 1.684560000000e-05, + 1.753370000000e-05, + 1.819940000000e-05, + 1.884250000000e-05, + 1.946310000000e-05,  \
+ 2.006150000000e-05, + 2.063790000000e-05, + 2.119280000000e-05, + 2.172660000000e-05, + 2.223980000000e-05,  \
+ 2.273290000000e-05, + 2.320660000000e-05, + 2.366140000000e-05, + 2.409810000000e-05, + 2.451710000000e-05,  \
+ 2.491930000000e-05, + 2.530510000000e-05, + 2.567520000000e-05, + 2.603040000000e-05, + 2.637100000000e-05,  \
+ 2.669790000000e-05, + 2.701140000000e-05, + 2.731220000000e-05, + 2.760090000000e-05, + 2.787790000000e-05,  \
+ 2.814370000000e-05, + 2.839880000000e-05, + 2.864380000000e-05, + 2.887890000000e-05, + 2.910460000000e-05,  \
+ 2.932140000000e-05, + 2.952950000000e-05, + 2.972950000000e-05, + 2.992160000000e-05, + 3.010610000000e-05 ]

.param id_pred_data_vd0.14=[ \
+ 3.116929470082e-10, + 4.488720684037e-10, + 6.508839778263e-10, + 9.466585915163e-10, + 1.378021270426e-09,  \
+ 2.006057293613e-09, + 2.920371890980e-09, + 4.251896967844e-09, + 6.190274035589e-09, + 9.007895442892e-09,  \
+ 1.309384259685e-08, + 1.900403105992e-08, + 2.753620350404e-08, + 3.983976114341e-08, + 5.756754319464e-08,  \
+ 8.306962399729e-08, + 1.196119274027e-07, + 1.715809662528e-07, + 2.446080361551e-07, + 3.455284740994e-07,  \
+ 4.821105585506e-07, + 6.625190872001e-07, + 8.945803529059e-07, + 1.184967077279e-06, + 1.538460728625e-06,  \
+ 1.957473814400e-06, + 2.441851247568e-06, + 2.989009772136e-06, + 3.594307345338e-06, + 4.251566970197e-06,  \
+ 4.953591997037e-06, + 5.692753111362e-06, + 6.461373632192e-06, + 7.252070499817e-06, + 8.058021412580e-06,  \
+ 8.873025944922e-06, + 9.691681771073e-06, + 1.050924052834e-05, + 1.132172546932e-05, + 1.212575574755e-05,  \
+ 1.291857595788e-05, + 1.369787787553e-05, + 1.446189722628e-05, + 1.520913458080e-05, + 1.593844397576e-05,  \
+ 1.664890762186e-05, + 1.733990007779e-05, + 1.801089674700e-05, + 1.866151054855e-05, + 1.929158868734e-05,  \
+ 1.990093151107e-05, + 2.048954309430e-05, + 2.105737454258e-05, + 2.160452364478e-05, + 2.213116560597e-05,  \
+ 2.263745933305e-05, + 2.312358206837e-05, + 2.358984347666e-05, + 2.403644524748e-05, + 2.446379279718e-05,  \
+ 2.487215708243e-05, + 2.526193333324e-05, + 2.563350659329e-05, + 2.598733728519e-05, + 2.632372692460e-05,  \
+ 2.664319297764e-05, + 2.694622846320e-05, + 2.723322249949e-05, + 2.750467217993e-05, + 2.776110923151e-05,  \
+ 2.800302667310e-05, + 2.823081362294e-05, + 2.844512404408e-05, + 2.864633075660e-05, + 2.883498789743e-05,  \
+ 2.901163126808e-05, + 2.917663776316e-05, + 2.933063689852e-05, + 2.947400556877e-05, + 2.960725920275e-05 ]

* Data table for Id-Vg at Vd = 0.15V
.param vg_data_vd0.15=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.15=[ \
+ 3.100540000000e-10, + 4.518770000000e-10, + 6.585570000000e-10, + 9.597330000000e-10, + 1.398600000000e-09,  \
+ 2.037900000000e-09, + 2.969200000000e-09, + 4.325400000000e-09, + 6.299600000000e-09, + 9.171700000000e-09,  \
+ 1.334680000000e-08, + 1.940880000000e-08, + 2.819520000000e-08, + 4.089960000000e-08, + 5.920510000000e-08,  \
+ 8.545220000000e-08, + 1.228330000000e-07, + 1.755820000000e-07, + 2.491240000000e-07, + 3.500790000000e-07,  \
+ 4.860710000000e-07, + 6.652510000000e-07, + 8.956010000000e-07, + 1.184100000000e-06, + 1.536100000000e-06,  \
+ 1.954800000000e-06, + 2.440800000000e-06, + 2.992700000000e-06, + 3.607000000000e-06, + 4.278700000000e-06,  \
+ 5.001500000000e-06, + 5.768500000000e-06, + 6.572200000000e-06, + 7.404900000000e-06, + 8.259300000000e-06,  \
+ 9.128100000000e-06, + 1.000470000000e-05, + 1.088290000000e-05, + 1.175750000000e-05, + 1.262380000000e-05,  \
+ 1.347810000000e-05, + 1.431720000000e-05, + 1.513860000000e-05, + 1.594060000000e-05, + 1.672180000000e-05,  \
+ 1.748120000000e-05, + 1.821810000000e-05, + 1.893220000000e-05, + 1.962320000000e-05, + 2.029110000000e-05,  \
+ 2.093610000000e-05, + 2.155830000000e-05, + 2.215800000000e-05, + 2.273560000000e-05, + 2.329160000000e-05,  \
+ 2.382650000000e-05, + 2.434070000000e-05, + 2.483500000000e-05, + 2.530990000000e-05, + 2.576600000000e-05,  \
+ 2.620390000000e-05, + 2.662440000000e-05, + 2.702790000000e-05, + 2.741530000000e-05, + 2.778700000000e-05,  \
+ 2.814380000000e-05, + 2.848620000000e-05, + 2.881470000000e-05, + 2.913000000000e-05, + 2.943260000000e-05,  \
+ 2.972300000000e-05, + 3.000180000000e-05, + 3.026940000000e-05, + 3.052620000000e-05, + 3.077290000000e-05,  \
+ 3.100960000000e-05, + 3.123700000000e-05, + 3.145540000000e-05, + 3.166510000000e-05, + 3.186650000000e-05 ]

.param id_pred_data_vd0.15=[ \
+ 3.164855377769e-10, + 4.555236521320e-10, + 6.602947522083e-10, + 9.600418460209e-10, + 1.397039151030e-09,  \
+ 2.033098622789e-09, + 2.959027156635e-09, + 4.307617729182e-09, + 6.271229935351e-09, + 9.125821165412e-09,  \
+ 1.326480365549e-08, + 1.924907380157e-08, + 2.788211688198e-08, + 4.031965374907e-08, + 5.822304132153e-08,  \
+ 8.395375061809e-08, + 1.207944080761e-07, + 1.731582642606e-07, + 2.467156889452e-07, + 3.483657906145e-07,  \
+ 4.859697924076e-07, + 6.678313411612e-07, + 9.019683602673e-07, + 1.195294589706e-06, + 1.552899539092e-06,  \
+ 1.977528609132e-06, + 2.469389710313e-06, + 3.026255035365e-06, + 3.643800482678e-06, + 4.316111790104e-06,  \
+ 5.036199945607e-06, + 5.796542245662e-06, + 6.589511758648e-06, + 7.407664088532e-06, + 8.244065065810e-06,  \
+ 9.092390064325e-06, + 9.946962745744e-06, + 1.080284673662e-05, + 1.165576977655e-05, + 1.250209643331e-05,  \
+ 1.333876862191e-05, + 1.416324666934e-05, + 1.497341436334e-05, + 1.576754839334e-05, + 1.654430634517e-05,  \
+ 1.730248986860e-05, + 1.804132953112e-05, + 1.876003298094e-05, + 1.945812764461e-05, + 2.013519770117e-05,  \
+ 2.079102487187e-05, + 2.142538432963e-05, + 2.203820622526e-05, + 2.262947964482e-05, + 2.319924169569e-05,  \
+ 2.374762771069e-05, + 2.427480794722e-05, + 2.478086753399e-05, + 2.526622774894e-05, + 2.573106758064e-05,  \
+ 2.617575810291e-05, + 2.660059835762e-05, + 2.700599652599e-05, + 2.739235424087e-05, + 2.776011024253e-05,  \
+ 2.810971418512e-05, + 2.844165937859e-05, + 2.875634309021e-05, + 2.905433284468e-05, + 2.933612631750e-05,  \
+ 2.960224301205e-05, + 2.985322862514e-05, + 3.008955027326e-05, + 3.031175365322e-05, + 3.052043030038e-05,  \
+ 3.071603860008e-05, + 3.089910678682e-05, + 3.107019801973e-05, + 3.122981215711e-05, + 3.137842504657e-05 ]

* Data table for Id-Vg at Vd = 0.16V
.param vg_data_vd0.16=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.16=[ \
+ 3.140550000000e-10, + 4.576570000000e-10, + 6.669050000000e-10, + 9.717900000000e-10, + 1.416000000000e-09,  \
+ 2.063100000000e-09, + 3.005500000000e-09, + 4.377800000000e-09, + 6.375100000000e-09, + 9.280600000000e-09,  \
+ 1.350370000000e-08, + 1.963450000000e-08, + 2.851970000000e-08, + 4.136520000000e-08, + 5.987130000000e-08,  \
+ 8.640230000000e-08, + 1.241810000000e-07, + 1.774840000000e-07, + 2.517840000000e-07, + 3.537650000000e-07,  \
+ 4.911180000000e-07, + 6.720740000000e-07, + 9.047000000000e-07, + 1.196100000000e-06, + 1.551700000000e-06,  \
+ 1.974800000000e-06, + 2.466200000000e-06, + 3.024800000000e-06, + 3.647200000000e-06, + 4.328800000000e-06,  \
+ 5.063600000000e-06, + 5.844900000000e-06, + 6.665700000000e-06, + 7.518600000000e-06, + 8.396400000000e-06,  \
+ 9.292000000000e-06, + 1.019890000000e-05, + 1.111080000000e-05, + 1.202210000000e-05, + 1.292790000000e-05,  \
+ 1.382390000000e-05, + 1.470670000000e-05, + 1.557320000000e-05, + 1.642140000000e-05, + 1.724930000000e-05,  \
+ 1.805570000000e-05, + 1.883970000000e-05, + 1.960080000000e-05, + 2.033850000000e-05, + 2.105260000000e-05,  \
+ 2.174320000000e-05, + 2.241030000000e-05, + 2.305420000000e-05, + 2.367520000000e-05, + 2.427360000000e-05,  \
+ 2.485000000000e-05, + 2.540480000000e-05, + 2.593850000000e-05, + 2.645170000000e-05, + 2.694500000000e-05,  \
+ 2.741900000000e-05, + 2.787440000000e-05, + 2.831180000000e-05, + 2.873180000000e-05, + 2.913510000000e-05,  \
+ 2.952230000000e-05, + 2.989390000000e-05, + 3.025070000000e-05, + 3.059320000000e-05, + 3.092190000000e-05,  \
+ 3.123740000000e-05, + 3.154030000000e-05, + 3.183100000000e-05, + 3.211020000000e-05, + 3.237810000000e-05,  \
+ 3.263540000000e-05, + 3.288240000000e-05, + 3.311950000000e-05, + 3.334730000000e-05, + 3.356600000000e-05 ]

.param id_pred_data_vd0.16=[ \
+ 3.210287857769e-10, + 4.618654614319e-10, + 6.693264964497e-10, + 9.729694028238e-10, + 1.415505579416e-09,  \
+ 2.059469892401e-09, + 2.996842454195e-09, + 4.362318293261e-09, + 6.350998660309e-09, + 9.242517080565e-09,  \
+ 1.343486133010e-08, + 1.949415946001e-08, + 2.822974238370e-08, + 4.080428880116e-08, + 5.888731266168e-08,  \
+ 8.485144462611e-08, + 1.219947716891e-07, + 1.747517853801e-07, + 2.488254176569e-07, + 3.511621980579e-07,  \
+ 4.896970131085e-07, + 6.728385051247e-07, + 9.087518265005e-07, + 1.204558648169e-06, + 1.565590500832e-06,  \
+ 1.994895574171e-06, + 2.493001229595e-06, + 3.058001166210e-06, + 3.685896517709e-06, + 4.371028626338e-06,  \
+ 5.106644821353e-06, + 5.885363207199e-06, + 6.699620280415e-06, + 7.542030652985e-06, + 8.405562839471e-06,  \
+ 9.283786057495e-06, + 1.017087721266e-05, + 1.106171403080e-05, + 1.195178483613e-05, + 1.283719786443e-05,  \
+ 1.371465972625e-05, + 1.458141021430e-05, + 1.543503371067e-05, + 1.627361285500e-05, + 1.709552132525e-05,  \
+ 1.789942034520e-05, + 1.868421211839e-05, + 1.944901072420e-05, + 2.019316656515e-05, + 2.091606846079e-05,  \
+ 2.161731943488e-05, + 2.229661447927e-05, + 2.295378362760e-05, + 2.358866855502e-05, + 2.420124597847e-05,  \
+ 2.479154150933e-05, + 2.535963896662e-05, + 2.590570133179e-05, + 2.642992418259e-05, + 2.693257993087e-05,  \
+ 2.741387579590e-05, + 2.787424949929e-05, + 2.831396181136e-05, + 2.873346908018e-05, + 2.913320204243e-05,  \
+ 2.951360540465e-05, + 2.987511688843e-05, + 3.021828364581e-05, + 3.054356435314e-05, + 3.085151081905e-05,  \
+ 3.114268649369e-05, + 3.141763852909e-05, + 3.167682560161e-05, + 3.192088566720e-05, + 3.215041942894e-05,  \
+ 3.236585529521e-05, + 3.256785683334e-05, + 3.275693161413e-05, + 3.293356625363e-05, + 3.309839870781e-05 ]

* Data table for Id-Vg at Vd = 0.17V
.param vg_data_vd0.17=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.17=[ \
+ 3.179690000000e-10, + 4.633080000000e-10, + 6.750620000000e-10, + 9.835630000000e-10, + 1.433000000000e-09,  \
+ 2.087600000000e-09, + 3.040900000000e-09, + 4.428800000000e-09, + 6.448600000000e-09, + 9.386500000000e-09,  \
+ 1.365610000000e-08, + 1.985370000000e-08, + 2.883450000000e-08, + 4.181630000000e-08, + 6.051620000000e-08,  \
+ 8.732070000000e-08, + 1.254820000000e-07, + 1.793160000000e-07, + 2.543410000000e-07, + 3.572970000000e-07,  \
+ 4.959370000000e-07, + 6.785600000000e-07, + 9.133040000000e-07, + 1.207400000000e-06, + 1.566200000000e-06,  \
+ 1.993300000000e-06, + 2.489600000000e-06, + 3.054000000000e-06, + 3.683500000000e-06, + 4.373600000000e-06,  \
+ 5.118600000000e-06, + 5.912100000000e-06, + 6.747400000000e-06, + 7.617400000000e-06, + 8.515200000000e-06,  \
+ 9.434000000000e-06, + 1.036700000000e-05, + 1.130830000000e-05, + 1.225220000000e-05, + 1.319330000000e-05,  \
+ 1.412730000000e-05, + 1.505020000000e-05, + 1.595870000000e-05, + 1.685020000000e-05, + 1.772240000000e-05,  \
+ 1.857370000000e-05, + 1.940300000000e-05, + 2.020940000000e-05, + 2.099230000000e-05, + 2.175140000000e-05,  \
+ 2.248650000000e-05, + 2.319760000000e-05, + 2.388490000000e-05, + 2.454860000000e-05, + 2.518890000000e-05,  \
+ 2.580630000000e-05, + 2.640120000000e-05, + 2.697420000000e-05, + 2.752560000000e-05, + 2.805610000000e-05,  \
+ 2.856630000000e-05, + 2.905690000000e-05, + 2.952830000000e-05, + 2.998120000000e-05, + 3.041630000000e-05,  \
+ 3.083430000000e-05, + 3.123560000000e-05, + 3.162100000000e-05, + 3.199100000000e-05, + 3.234630000000e-05,  \
+ 3.268730000000e-05, + 3.301480000000e-05, + 3.332910000000e-05, + 3.363090000000e-05, + 3.392060000000e-05,  \
+ 3.419870000000e-05, + 3.446570000000e-05, + 3.472200000000e-05, + 3.496810000000e-05, + 3.520440000000e-05 ]

.param id_pred_data_vd0.17=[ \
+ 3.253566083217e-10, + 4.679365894766e-10, + 6.780302364007e-10, + 9.855070226550e-10, + 1.433510510296e-09,  \
+ 2.085275978558e-09, + 3.033966198274e-09, + 4.416163097432e-09, + 6.429819379150e-09, + 9.358365637979e-09,  \
+ 1.360450426091e-08, + 1.973997584059e-08, + 2.858047665200e-08, + 4.129592809932e-08, + 5.956484017133e-08,  \
+ 8.577091534789e-08, + 1.232270409446e-07, + 1.763870307059e-07, + 2.509804676265e-07, + 3.539911836015e-07,  \
+ 4.934076446261e-07, + 6.777203680031e-07, + 9.152091706710e-07, + 1.213151390402e-06, + 1.577091024956e-06,  \
+ 2.010320349655e-06, + 2.513655417715e-06, + 3.085495354753e-06, + 3.722119527083e-06, + 4.418149837875e-06,  \
+ 5.167064664420e-06, + 5.961656206637e-06, + 6.794479486416e-06, + 7.658189097128e-06, + 8.545771743229e-06,  \
+ 9.450705183554e-06, + 1.036706460582e-05, + 1.128956653702e-05, + 1.221354657901e-05, + 1.313490189204e-05,  \
+ 1.405013324984e-05, + 1.495618918852e-05, + 1.585054640600e-05, + 1.673096361628e-05, + 1.759562626830e-05,  \
+ 1.844299564254e-05, + 1.927175318997e-05, + 2.008087103604e-05, + 2.086943510221e-05, + 2.163675890188e-05,  \
+ 2.238222645246e-05, + 2.310542462510e-05, + 2.380606398219e-05, + 2.448387240293e-05, + 2.513872372219e-05,  \
+ 2.577055856818e-05, + 2.637937446707e-05, + 2.696526047657e-05, + 2.752837739536e-05, + 2.806883654557e-05,  \
+ 2.858703621314e-05, + 2.908316688263e-05, + 2.955767384265e-05, + 3.001079952810e-05, + 3.044296201551e-05,  \
+ 3.085470554652e-05, + 3.124649767415e-05, + 3.161877131788e-05, + 3.197205587639e-05, + 3.230691043427e-05,  \
+ 3.262385944254e-05, + 3.292350156698e-05, + 3.320641568280e-05, + 3.347314603161e-05, + 3.372425911948e-05,  \
+ 3.396044514375e-05, + 3.418210981181e-05, + 3.439000269282e-05, + 3.458457649685e-05, + 3.476648926153e-05 ]

* Data table for Id-Vg at Vd = 0.18V
.param vg_data_vd0.18=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.18=[ \
+ 3.218200000000e-10, + 4.688650000000e-10, + 6.830790000000e-10, + 9.951280000000e-10, + 1.449700000000e-09,  \
+ 2.111600000000e-09, + 3.075500000000e-09, + 4.478700000000e-09, + 6.520600000000e-09, + 9.490100000000e-09,  \
+ 1.380520000000e-08, + 2.006800000000e-08, + 2.914200000000e-08, + 4.225660000000e-08, + 6.114490000000e-08,  \
+ 8.821510000000e-08, + 1.267480000000e-07, + 1.810940000000e-07, + 2.568180000000e-07, + 3.607100000000e-07,  \
+ 5.005790000000e-07, + 6.847830000000e-07, + 9.215230000000e-07, + 1.218000000000e-06, + 1.579900000000e-06,  \
+ 2.010600000000e-06, + 2.511300000000e-06, + 3.080900000000e-06, + 3.716700000000e-06, + 4.414200000000e-06,  \
+ 5.168100000000e-06, + 5.972100000000e-06, + 6.819900000000e-06, + 7.704600000000e-06, + 8.619500000000e-06,  \
+ 9.558000000000e-06, + 1.051380000000e-05, + 1.148070000000e-05, + 1.245310000000e-05, + 1.342570000000e-05,  \
+ 1.439380000000e-05, + 1.535320000000e-05, + 1.630030000000e-05, + 1.723200000000e-05, + 1.814580000000e-05,  \
+ 1.903980000000e-05, + 1.991230000000e-05, + 2.076220000000e-05, + 2.158880000000e-05, + 2.239140000000e-05,  \
+ 2.316980000000e-05, + 2.392390000000e-05, + 2.465360000000e-05, + 2.535910000000e-05, + 2.604060000000e-05,  \
+ 2.669850000000e-05, + 2.733300000000e-05, + 2.794480000000e-05, + 2.853420000000e-05, + 2.910170000000e-05,  \
+ 2.964800000000e-05, + 3.017360000000e-05, + 3.067910000000e-05, + 3.116500000000e-05, + 3.163220000000e-05,  \
+ 3.208110000000e-05, + 3.251230000000e-05, + 3.292660000000e-05, + 3.332450000000e-05, + 3.370660000000e-05,  \
+ 3.407350000000e-05, + 3.442590000000e-05, + 3.476410000000e-05, + 3.508890000000e-05, + 3.540060000000e-05,  \
+ 3.569990000000e-05, + 3.598730000000e-05, + 3.626310000000e-05, + 3.652780000000e-05, + 3.678200000000e-05 ]

.param id_pred_data_vd0.18=[ \
+ 3.294980288615e-10, + 4.737681447153e-10, + 6.864421031594e-10, + 9.976935277933e-10, + 1.451093005755e-09,  \
+ 2.110558767754e-09, + 3.070429031027e-09, + 4.469186620781e-09, + 6.507665446520e-09, + 9.473222206680e-09,  \
+ 1.377352248255e-08, + 1.998634346023e-08, + 2.893406218618e-08, + 4.179474558441e-08, + 6.025651146047e-08,  \
+ 8.671494242662e-08, + 1.244976908765e-07, + 1.780772367965e-07, + 2.532054872972e-07, + 3.568958300093e-07,  \
+ 4.971783573637e-07, + 6.826000935689e-07, + 9.215299269272e-07, + 1.221366810569e-06, + 1.587817969266e-06,  \
+ 2.024387595156e-06, + 2.532133494242e-06, + 3.109730605502e-06, + 3.753720739041e-06, + 4.459014344320e-06,  \
+ 5.219289305387e-06, + 6.027547715348e-06, + 6.876484549139e-06, + 7.758820647723e-06, + 8.667600341141e-06,  \
+ 9.596263480489e-06, + 1.053885105648e-05, + 1.148991286755e-05, + 1.244468890945e-05, + 1.339890834060e-05,  \
+ 1.434887919459e-05, + 1.529136919999e-05, + 1.622359923203e-05, + 1.714321842883e-05, + 1.804814441130e-05,  \
+ 1.893665496027e-05, + 1.980723085580e-05, + 2.065864100587e-05, + 2.148984553060e-05, + 2.229998266557e-05,  \
+ 2.308830851689e-05, + 2.385415253229e-05, + 2.459718991304e-05, + 2.531704871217e-05, + 2.601343032438e-05,  \
+ 2.668622735655e-05, + 2.733530884143e-05, + 2.796073764330e-05, + 2.856256352970e-05, + 2.914091222920e-05,  \
+ 2.969600376673e-05, + 3.022809483809e-05, + 3.073751810007e-05, + 3.122457215795e-05, + 3.168968134560e-05,  \
+ 3.213320713257e-05, + 3.255569958128e-05, + 3.295767994132e-05, + 3.333955944981e-05, + 3.370200865902e-05,  \
+ 3.404546761885e-05, + 3.437058854615e-05, + 3.467790840659e-05, + 3.496806108160e-05, + 3.524161234964e-05,  \
+ 3.549922228558e-05, + 3.574146190658e-05, + 3.596892056521e-05, + 3.618215880124e-05, + 3.638191003120e-05 ]

* Data table for Id-Vg at Vd = 0.19V
.param vg_data_vd0.19=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.19=[ \
+ 3.256270000000e-10, + 4.743550000000e-10, + 6.909970000000e-10, + 1.006500000000e-09, + 1.466100000000e-09,  \
+ 2.135300000000e-09, + 3.109700000000e-09, + 4.528000000000e-09, + 6.591500000000e-09, + 9.592100000000e-09,  \
+ 1.395180000000e-08, + 2.027850000000e-08, + 2.944390000000e-08, + 4.268860000000e-08, + 6.176120000000e-08,  \
+ 8.909080000000e-08, + 1.279860000000e-07, + 1.828310000000e-07, + 2.592330000000e-07, + 3.640290000000e-07,  \
+ 5.050810000000e-07, + 6.907990000000e-07, + 9.294350000000e-07, + 1.228300000000e-06, + 1.593000000000e-06,  \
+ 2.027100000000e-06, + 2.531700000000e-06, + 3.106100000000e-06, + 3.747400000000e-06, + 4.451500000000e-06,  \
+ 5.213200000000e-06, + 6.026400000000e-06, + 6.884900000000e-06, + 7.782300000000e-06, + 8.711900000000e-06,  \
+ 9.667600000000e-06, + 1.064290000000e-05, + 1.163210000000e-05, + 1.262960000000e-05, + 1.362990000000e-05,  \
+ 1.462850000000e-05, + 1.562080000000e-05, + 1.660310000000e-05, + 1.757190000000e-05, + 1.852440000000e-05,  \
+ 1.945830000000e-05, + 2.037180000000e-05, + 2.126330000000e-05, + 2.213170000000e-05, + 2.297640000000e-05,  \
+ 2.379680000000e-05, + 2.459260000000e-05, + 2.536360000000e-05, + 2.611000000000e-05, + 2.683190000000e-05,  \
+ 2.752950000000e-05, + 2.820320000000e-05, + 2.885320000000e-05, + 2.948010000000e-05, + 3.008430000000e-05,  \
+ 3.066640000000e-05, + 3.122680000000e-05, + 3.176630000000e-05, + 3.228520000000e-05, + 3.278440000000e-05,  \
+ 3.326430000000e-05, + 3.372560000000e-05, + 3.416890000000e-05, + 3.459490000000e-05, + 3.500410000000e-05,  \
+ 3.539710000000e-05, + 3.577450000000e-05, + 3.613700000000e-05, + 3.648500000000e-05, + 3.681910000000e-05,  \
+ 3.713980000000e-05, + 3.744770000000e-05, + 3.774330000000e-05, + 3.802700000000e-05, + 3.829920000000e-05 ]

.param id_pred_data_vd0.19=[ \
+ 3.334754039575e-10, + 4.793900876265e-10, + 6.945916841694e-10, + 1.009561514387e-09, + 1.468289880791e-09,  \
+ 2.135355146038e-09, + 3.106259782726e-09, + 4.521391847589e-09, + 6.584486236250e-09, + 9.586969795805e-09,  \
+ 1.394167092883e-08, + 2.023265295747e-08, + 2.928972065774e-08, + 4.229965540503e-08, + 6.096107455278e-08,  \
+ 8.768253906055e-08, + 1.258070636823e-07, + 1.798253975949e-07, + 2.555107926128e-07, + 3.599000649501e-07,  \
+ 5.010527388549e-07, + 6.875586632304e-07, + 9.278471088692e-07, + 1.229409863299e-06, + 1.598083727004e-06,  \
+ 2.037540180027e-06, + 2.549044147599e-06, + 3.131511111860e-06, + 3.781742470892e-06, + 4.494872064242e-06,  \
+ 5.264839655865e-06, + 6.084828128223e-06, + 6.947693764232e-06, + 7.846264161344e-06, + 8.773649278737e-06,  \
+ 9.723323346407e-06, + 1.068925204891e-05, + 1.166595196992e-05, + 1.264854588953e-05, + 1.363266324915e-05,  \
+ 1.461441941501e-05, + 1.559047443152e-05, + 1.655781183217e-05, + 1.751393770974e-05, + 1.845657105150e-05,  \
+ 1.938377645274e-05, + 2.029392402619e-05, + 2.118558018992e-05, + 2.205749937275e-05, + 2.290866963449e-05,  \
+ 2.373817857006e-05, + 2.454537228914e-05, + 2.532957340009e-05, + 2.609036440845e-05, + 2.682742735487e-05,  \
+ 2.754039174761e-05, + 2.822916911100e-05, + 2.889364332077e-05, + 2.953385032015e-05, + 3.014980393345e-05,  \
+ 3.074172811466e-05, + 3.130975004751e-05, + 3.185422639945e-05, + 3.237539771362e-05, + 3.287366489531e-05,  \
+ 3.334937355248e-05, + 3.380306836334e-05, + 3.423517235206e-05, + 3.464619425358e-05, + 3.503677828121e-05,  \
+ 3.540734469425e-05, + 3.575856258976e-05, + 3.609102641349e-05, + 3.640525595983e-05, + 3.670205303933e-05,  \
+ 3.698183514643e-05, + 3.724527137820e-05, + 3.749313313165e-05, + 3.772591255256e-05, + 3.794424555963e-05 ]

* Data table for Id-Vg at Vd = 0.20V
.param vg_data_vd0.20=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.20=[ \
+ 3.294040000000e-10, + 4.797990000000e-10, + 6.988440000000e-10, + 1.017900000000e-09, + 1.482400000000e-09,  \
+ 2.158800000000e-09, + 3.143500000000e-09, + 4.576600000000e-09, + 6.661500000000e-09, + 9.692800000000e-09,  \
+ 1.409650000000e-08, + 2.048620000000e-08, + 2.974150000000e-08, + 4.311420000000e-08, + 6.236790000000e-08,  \
+ 8.995210000000e-08, + 1.292020000000e-07, + 1.845350000000e-07, + 2.615980000000e-07, + 3.672730000000e-07,  \
+ 5.094710000000e-07, + 6.966480000000e-07, + 9.371010000000e-07, + 1.238200000000e-06, + 1.605500000000e-06,  \
+ 2.042800000000e-06, + 2.551100000000e-06, + 3.129800000000e-06, + 3.776200000000e-06, + 4.486200000000e-06,  \
+ 5.254800000000e-06, + 6.076100000000e-06, + 6.944000000000e-06, + 7.852400000000e-06, + 8.794900000000e-06,  \
+ 9.765300000000e-06, + 1.075770000000e-05, + 1.176630000000e-05, + 1.278560000000e-05, + 1.381050000000e-05,  \
+ 1.483600000000e-05, + 1.585780000000e-05, + 1.687190000000e-05, + 1.787460000000e-05, + 1.886280000000e-05,  \
+ 1.983400000000e-05, + 2.078590000000e-05, + 2.171670000000e-05, + 2.262520000000e-05, + 2.351020000000e-05,  \
+ 2.437100000000e-05, + 2.520720000000e-05, + 2.601850000000e-05, + 2.680480000000e-05, + 2.756610000000e-05,  \
+ 2.830270000000e-05, + 2.901460000000e-05, + 2.970230000000e-05, + 3.036620000000e-05, + 3.100660000000e-05,  \
+ 3.162400000000e-05, + 3.221900000000e-05, + 3.279220000000e-05, + 3.334400000000e-05, + 3.387500000000e-05,  \
+ 3.438590000000e-05, + 3.487720000000e-05, + 3.534960000000e-05, + 3.580370000000e-05, + 3.624010000000e-05,  \
+ 3.665930000000e-05, + 3.706200000000e-05, + 3.744880000000e-05, + 3.782030000000e-05, + 3.817690000000e-05,  \
+ 3.851930000000e-05, + 3.884800000000e-05, + 3.916350000000e-05, + 3.946620000000e-05, + 3.975680000000e-05 ]

.param id_pred_data_vd0.20=[ \
+ 3.373139323415e-10, + 4.848259127499e-10, + 7.025065418276e-10, + 1.021143258839e-09, + 1.485128553469e-09,  \
+ 2.159691447901e-09, + 3.141463622569e-09, + 4.572720868623e-09, + 6.660125961844e-09, + 9.699265035579e-09,  \
+ 1.410836460991e-08, + 2.047804059657e-08, + 2.964603140754e-08, + 4.280855421257e-08, + 6.167583705974e-08,  \
+ 8.867025940162e-08, + 1.271517135137e-07, + 1.816297526602e-07, + 2.578971816547e-07, + 3.630113724284e-07,  \
+ 5.050542768004e-07, + 6.926426522114e-07, + 9.342479643237e-07, + 1.237423748535e-06, + 1.608106504136e-06,  \
+ 2.050108014373e-06, + 2.564862552390e-06, + 3.151478813379e-06, + 3.807003304246e-06, + 4.526795964921e-06,  \
+ 5.305013837642e-06, + 6.135043076938e-06, + 7.009915134404e-06, + 7.922582881292e-06, + 8.866240386851e-06,  \
+ 9.834392403718e-06, + 1.082103044610e-05, + 1.182064443128e-05, + 1.282826415263e-05, + 1.383943745168e-05,  \
+ 1.485015527578e-05, + 1.585691788932e-05, + 1.685663009994e-05, + 1.784656342352e-05, + 1.882430806290e-05,  \
+ 1.978781365324e-05, + 2.073519572150e-05, + 2.166484919144e-05, + 2.257547312183e-05, + 2.346580149606e-05,  \
+ 2.433483023196e-05, + 2.518175751902e-05, + 2.600572770461e-05, + 2.680627512746e-05, + 2.758284099400e-05,  \
+ 2.833511098288e-05, + 2.906274457928e-05, + 2.976565447170e-05, + 3.044375916943e-05, + 3.109695098829e-05,  \
+ 3.172537835781e-05, + 3.232926828787e-05, + 3.290873137303e-05, + 3.346406447235e-05, + 3.399558481760e-05,  \
+ 3.450371441431e-05, + 3.498892474454e-05, + 3.545157087501e-05, + 3.589218249545e-05, + 3.631132130977e-05,  \
+ 3.670950827654e-05, + 3.708743606694e-05, + 3.744560526684e-05, + 3.778467071243e-05, + 3.810521448031e-05,  \
+ 3.840795834549e-05, + 3.869343781844e-05, + 3.896234265994e-05, + 3.921538300347e-05, + 3.945305943489e-05 ]

* Data table for Id-Vg at Vd = 0.21V
.param vg_data_vd0.21=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.21=[ \
+ 3.331600000000e-10, + 4.852120000000e-10, + 7.066430000000e-10, + 1.029100000000e-09, + 1.498600000000e-09,  \
+ 2.182100000000e-09, + 3.177100000000e-09, + 4.624900000000e-09, + 6.730900000000e-09, + 9.792600000000e-09,  \
+ 1.423980000000e-08, + 2.069180000000e-08, + 3.003590000000e-08, + 4.353490000000e-08, + 6.296720000000e-08,  \
+ 9.080210000000e-08, + 1.304000000000e-07, + 1.862120000000e-07, + 2.639230000000e-07, + 3.704580000000e-07,  \
+ 5.137700000000e-07, + 7.023610000000e-07, + 9.445670000000e-07, + 1.247800000000e-06, + 1.617700000000e-06,  \
+ 2.057800000000e-06, + 2.569700000000e-06, + 3.152400000000e-06, + 3.803400000000e-06, + 4.518800000000e-06,  \
+ 5.293500000000e-06, + 6.122000000000e-06, + 6.998300000000e-06, + 7.916400000000e-06, + 8.870100000000e-06,  \
+ 9.853400000000e-06, + 1.086070000000e-05, + 1.188630000000e-05, + 1.292480000000e-05, + 1.397110000000e-05,  \
+ 1.502060000000e-05, + 1.606860000000e-05, + 1.711120000000e-05, + 1.814470000000e-05, + 1.916560000000e-05,  \
+ 2.017110000000e-05, + 2.115880000000e-05, + 2.212670000000e-05, + 2.307300000000e-05, + 2.399650000000e-05,  \
+ 2.489610000000e-05, + 2.577130000000e-05, + 2.662160000000e-05, + 2.744660000000e-05, + 2.824640000000e-05,  \
+ 2.902090000000e-05, + 2.977040000000e-05, + 3.049510000000e-05, + 3.119520000000e-05, + 3.187130000000e-05,  \
+ 3.252360000000e-05, + 3.315280000000e-05, + 3.375920000000e-05, + 3.434350000000e-05, + 3.490620000000e-05,  \
+ 3.544790000000e-05, + 3.596920000000e-05, + 3.647060000000e-05, + 3.695270000000e-05, + 3.741630000000e-05,  \
+ 3.786180000000e-05, + 3.828980000000e-05, + 3.870110000000e-05, + 3.909600000000e-05, + 3.947530000000e-05,  \
+ 3.983950000000e-05, + 4.018910000000e-05, + 4.052460000000e-05, + 4.084660000000e-05, + 4.115560000000e-05 ]

.param id_pred_data_vd0.21=[ \
+ 3.410337612308e-10, + 4.901032779614e-10, + 7.102143606552e-10, + 1.032465299922e-09, + 1.501638053902e-09,  \
+ 2.183587231031e-09, + 3.176034368835e-09, + 4.623148051053e-09, + 6.734497439709e-09, + 9.809836996055e-09,  \
+ 1.427298364831e-08, + 2.072140880216e-08, + 3.000138846687e-08, + 4.331908186828e-08, + 6.239714792855e-08,  \
+ 8.967357587153e-08, + 1.285259702399e-07, + 1.834830646885e-07, + 2.603583311611e-07, + 3.662275798888e-07,  \
+ 5.091874118079e-07, + 6.978735677876e-07, + 9.407794505023e-07, + 1.245505613952e-06, + 1.618053802304e-06,  \
+ 2.062333087451e-06, + 2.579935498943e-06, + 3.170138315909e-06, + 3.830179957731e-06, + 4.555631276162e-06,  \
+ 5.340884308680e-06, + 6.179495685501e-06, + 7.064686651574e-06, + 7.989558507688e-06, + 8.947377573350e-06,  \
+ 9.931756248989e-06, + 1.093669045076e-05, + 1.195667726279e-05, + 1.298668743402e-05, + 1.402221962053e-05,  \
+ 1.505920488853e-05, + 1.609399449080e-05, + 1.712339348160e-05, + 1.814450792153e-05, + 1.915480905154e-05,  \
+ 2.015209662204e-05, + 2.113436748914e-05, + 2.209982325439e-05, + 2.304701083631e-05, + 2.397453979938e-05,  \
+ 2.488124278898e-05, + 2.576617553132e-05, + 2.662843500730e-05, + 2.746729238424e-05, + 2.828220371157e-05,  \
+ 2.907264643000e-05, + 2.983824771945e-05, + 3.057868976612e-05, + 3.129399396130e-05, + 3.198390666512e-05,  \
+ 3.264846760430e-05, + 3.328779595904e-05, + 3.390215453692e-05, + 3.449158000876e-05, + 3.505640241201e-05,  \
+ 3.559704957297e-05, + 3.611389125581e-05, + 3.660729111289e-05, + 3.707785726874e-05, + 3.752601143788e-05,  \
+ 3.795228229137e-05, + 3.835737879854e-05, + 3.874177768012e-05, + 3.910619096132e-05, + 3.945114731323e-05,  \
+ 3.977744432632e-05, + 4.008556177723e-05, + 4.037626975332e-05, + 4.065020082635e-05, + 4.090799979167e-05 ]

* Data table for Id-Vg at Vd = 0.22V
.param vg_data_vd0.22=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.22=[ \
+ 3.369040000000e-10, + 4.906050000000e-10, + 7.144110000000e-10, + 1.040300000000e-09, + 1.514700000000e-09,  \
+ 2.205300000000e-09, + 3.210400000000e-09, + 4.672900000000e-09, + 6.799900000000e-09, + 9.891700000000e-09,  \
+ 1.438210000000e-08, + 2.089580000000e-08, + 3.032790000000e-08, + 4.395180000000e-08, + 6.356070000000e-08,  \
+ 9.164320000000e-08, + 1.315850000000e-07, + 1.878690000000e-07, + 2.662170000000e-07, + 3.735940000000e-07,  \
+ 5.179960000000e-07, + 7.079640000000e-07, + 9.518670000000e-07, + 1.257100000000e-06, + 1.629400000000e-06,  \
+ 2.072400000000e-06, + 2.587500000000e-06, + 3.174000000000e-06, + 3.829300000000e-06, + 4.549600000000e-06,  \
+ 5.329900000000e-06, + 6.164900000000e-06, + 7.048700000000e-06, + 7.975300000000e-06, + 8.938900000000e-06,  \
+ 9.933700000000e-06, + 1.095400000000e-05, + 1.199440000000e-05, + 1.304970000000e-05, + 1.411510000000e-05,  \
+ 1.518570000000e-05, + 1.625710000000e-05, + 1.732530000000e-05, + 1.838640000000e-05, + 1.943700000000e-05,  \
+ 2.047410000000e-05, + 2.149490000000e-05, + 2.249720000000e-05, + 2.347910000000e-05, + 2.443900000000e-05,  \
+ 2.537580000000e-05, + 2.628830000000e-05, + 2.717610000000e-05, + 2.803870000000e-05, + 2.887580000000e-05,  \
+ 2.968740000000e-05, + 3.047350000000e-05, + 3.123430000000e-05, + 3.197010000000e-05, + 3.268110000000e-05,  \
+ 3.336780000000e-05, + 3.403060000000e-05, + 3.467000000000e-05, + 3.528640000000e-05, + 3.588050000000e-05,  \
+ 3.645260000000e-05, + 3.700360000000e-05, + 3.753380000000e-05, + 3.804390000000e-05, + 3.853450000000e-05,  \
+ 3.900620000000e-05, + 3.945960000000e-05, + 3.989520000000e-05, + 4.031380000000e-05, + 4.071580000000e-05,  \
+ 4.110180000000e-05, + 4.147230000000e-05, + 4.182800000000e-05, + 4.216930000000e-05, + 4.249680000000e-05 ]

.param id_pred_data_vd0.22=[ \
+ 3.446564122989e-10, + 4.952442411721e-10, + 7.177449301565e-10, + 1.043556085989e-09, + 1.517843903898e-09,  \
+ 2.207068749982e-09, + 3.210004457799e-09, + 4.672640940839e-09, + 6.807462966663e-09, + 9.918449634938e-09,  \
+ 1.443505723842e-08, + 2.096198315371e-08, + 3.035410145458e-08, + 4.382857440532e-08, + 6.312145558240e-08,  \
+ 9.068683141322e-08, + 1.299219695738e-07, + 1.853765900250e-07, + 2.628841889418e-07, + 3.695372902257e-07,  \
+ 5.134457569511e-07, + 7.032543271634e-07, + 9.474672515353e-07, + 1.253707914657e-06, + 1.628023101148e-06,  \
+ 2.074400581478e-06, + 2.594536908873e-06, + 3.187864131178e-06, + 3.851798101095e-06, + 4.582100336847e-06,  \
+ 5.373334824981e-06, + 6.219300812518e-06, + 7.113347746781e-06, + 8.048741437960e-06, + 9.018875352922e-06,  \
+ 1.001742268272e-05, + 1.103845519538e-05, + 1.207649846037e-05, + 1.312646621955e-05, + 1.418387968442e-05,  \
+ 1.524453458842e-05, + 1.630475890124e-05, + 1.736125836032e-05, + 1.841101882746e-05, + 1.945140233147e-05,  \
+ 2.048002381343e-05, + 2.149475432816e-05, + 2.249372104416e-05, + 2.347531364649e-05, + 2.443799545290e-05,  \
+ 2.538046988775e-05, + 2.630161165143e-05, + 2.720046031754e-05, + 2.807615790516e-05, + 2.892796648666e-05,  \
+ 2.975532261189e-05, + 3.055778128328e-05, + 3.133499034448e-05, + 3.208658163203e-05, + 3.281255194452e-05,  \
+ 3.351270279381e-05, + 3.418714302825e-05, + 3.483583423076e-05, + 3.545914136339e-05, + 3.605720208725e-05,  \
+ 3.663025971036e-05, + 3.717879764736e-05, + 3.770317445742e-05, + 3.820374869974e-05, + 3.868125990266e-05,  \
+ 3.913595457561e-05, + 3.956862346968e-05, + 3.997972438810e-05, + 4.036998405354e-05, + 4.073995951330e-05,  \
+ 4.109035508009e-05, + 4.142175341258e-05, + 4.173488443485e-05, + 4.203033720842e-05, + 4.230891208863e-05 ]

* Data table for Id-Vg at Vd = 0.23V
.param vg_data_vd0.23=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.23=[ \
+ 3.406420000000e-10, + 4.959880000000e-10, + 7.221610000000e-10, + 1.051400000000e-09, + 1.530700000000e-09,  \
+ 2.228400000000e-09, + 3.243600000000e-09, + 4.720600000000e-09, + 6.868600000000e-09, + 9.990300000000e-09,  \
+ 1.452360000000e-08, + 2.109860000000e-08, + 3.061800000000e-08, + 4.436590000000e-08, + 6.414970000000e-08,  \
+ 9.247740000000e-08, + 1.327600000000e-07, + 1.895100000000e-07, + 2.684840000000e-07, + 3.766900000000e-07,  \
+ 5.221620000000e-07, + 7.134750000000e-07, + 9.590310000000e-07, + 1.266300000000e-06, + 1.640900000000e-06,  \
+ 2.086600000000e-06, + 2.604800000000e-06, + 3.194800000000e-06, + 3.854100000000e-06, + 4.578900000000e-06,  \
+ 5.364500000000e-06, + 6.205300000000e-06, + 7.095800000000e-06, + 8.030100000000e-06, + 9.002500000000e-06,  \
+ 1.000730000000e-05, + 1.103920000000e-05, + 1.209270000000e-05, + 1.316290000000e-05, + 1.424500000000e-05,  \
+ 1.533430000000e-05, + 1.642650000000e-05, + 1.751750000000e-05, + 1.860350000000e-05, + 1.968100000000e-05,  \
+ 2.074680000000e-05, + 2.179810000000e-05, + 2.283240000000e-05, + 2.384750000000e-05, + 2.484170000000e-05,  \
+ 2.581340000000e-05, + 2.676160000000e-05, + 2.768540000000e-05, + 2.858420000000e-05, + 2.945740000000e-05,  \
+ 3.030500000000e-05, + 3.112680000000e-05, + 3.192300000000e-05, + 3.269360000000e-05, + 3.343890000000e-05,  \
+ 3.415930000000e-05, + 3.485520000000e-05, + 3.552700000000e-05, + 3.617510000000e-05, + 3.680000000000e-05,  \
+ 3.740240000000e-05, + 3.798260000000e-05, + 3.854140000000e-05, + 3.907920000000e-05, + 3.959680000000e-05,  \
+ 4.009450000000e-05, + 4.057310000000e-05, + 4.103310000000e-05, + 4.147510000000e-05, + 4.189980000000e-05,  \
+ 4.230760000000e-05, + 4.269910000000e-05, + 4.307490000000e-05, + 4.343560000000e-05, + 4.378160000000e-05 ]

.param id_pred_data_vd0.23=[ \
+ 3.482016996958e-10, + 5.002746061855e-10, + 7.251252620577e-10, + 1.054451521654e-09, + 1.533793603237e-09,  \
+ 2.230175706330e-09, + 3.243395347852e-09, + 4.721210125069e-09, + 6.878983320746e-09, + 1.002491046620e-08,  \
+ 1.459417227068e-08, + 2.119878573126e-08, + 3.070279916528e-08, + 4.433464269482e-08, + 6.384462892584e-08,  \
+ 9.170447015094e-08, + 1.313317750373e-07, + 1.872991833807e-07, + 2.654612262631e-07, + 3.729268053121e-07,  \
+ 5.178163564779e-07, + 7.087761514413e-07, + 9.543148189550e-07, + 1.262058467546e-06, + 1.638082421778e-06,  \
+ 2.086425811285e-06, + 2.608868371681e-06, + 3.204965378245e-06, + 3.872272936860e-06, + 4.606746897480e-06,  \
+ 5.403123777796e-06, + 6.255366115511e-06, + 7.157013060350e-06, + 8.101478670142e-06, + 9.082289543585e-06,  \
+ 1.009320865705e-05, + 1.112836380344e-05, + 1.218230616360e-05, + 1.325005130639e-05, + 1.432698045392e-05,  \
+ 1.540892750199e-05, + 1.649215642828e-05, + 1.757326339430e-05, + 1.864921439847e-05, + 1.971717290871e-05,  \
+ 2.077474418911e-05, + 2.181963558542e-05, + 2.284984395374e-05, + 2.386360712990e-05, + 2.485939388862e-05,  \
+ 2.583563116787e-05, + 2.679114753846e-05, + 2.772483014269e-05, + 2.863570000045e-05, + 2.952297727461e-05,  \
+ 3.038592229132e-05, + 3.122402296867e-05, + 3.203671367373e-05, + 3.282376012066e-05, + 3.358485104400e-05,  \
+ 3.431986930082e-05, + 3.502872452373e-05, + 3.571149703930e-05, + 3.636826048023e-05, + 3.699925917317e-05,  \
+ 3.760460691410e-05, + 3.818477227469e-05, + 3.874003639794e-05, + 3.927084777388e-05, + 3.977774191299e-05,  \
+ 4.026114052976e-05, + 4.072166615515e-05, + 4.115989111597e-05, + 4.157642120845e-05, + 4.197177855531e-05,  \
+ 4.234673964675e-05, + 4.270199395251e-05, + 4.303806024836e-05, + 4.335571837146e-05, + 4.365565109765e-05 ]

* Data table for Id-Vg at Vd = 0.24V
.param vg_data_vd0.24=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.24=[ \
+ 3.443790000000e-10, + 5.013680000000e-10, + 7.299040000000e-10, + 1.062600000000e-09, + 1.546800000000e-09,  \
+ 2.251500000000e-09, + 3.276800000000e-09, + 4.768300000000e-09, + 6.937000000000e-09, + 1.008860000000e-08,  \
+ 1.466460000000e-08, + 2.130050000000e-08, + 3.090670000000e-08, + 4.477780000000e-08, + 6.473530000000e-08,  \
+ 9.330630000000e-08, + 1.339260000000e-07, + 1.911370000000e-07, + 2.707310000000e-07, + 3.797540000000e-07,  \
+ 5.262770000000e-07, + 7.189090000000e-07, + 9.660790000000e-07, + 1.275200000000e-06, + 1.652100000000e-06,  \
+ 2.100500000000e-06, + 2.621600000000e-06, + 3.214900000000e-06, + 3.878000000000e-06, + 4.607100000000e-06,  \
+ 5.397400000000e-06, + 6.243600000000e-06, + 7.140200000000e-06, + 8.081400000000e-06, + 9.061800000000e-06,  \
+ 1.007560000000e-05, + 1.111770000000e-05, + 1.218290000000e-05, + 1.326620000000e-05, + 1.436310000000e-05,  \
+ 1.546900000000e-05, + 1.657970000000e-05, + 1.769110000000e-05, + 1.879950000000e-05, + 1.990120000000e-05,  \
+ 2.099310000000e-05, + 2.207220000000e-05, + 2.313590000000e-05, + 2.418180000000e-05, + 2.520800000000e-05,  \
+ 2.621280000000e-05, + 2.719470000000e-05, + 2.815280000000e-05, + 2.908620000000e-05, + 2.999430000000e-05,  \
+ 3.087670000000e-05, + 3.173320000000e-05, + 3.256370000000e-05, + 3.336830000000e-05, + 3.414720000000e-05,  \
+ 3.490070000000e-05, + 3.562900000000e-05, + 3.633260000000e-05, + 3.701190000000e-05, + 3.766730000000e-05,  \
+ 3.829940000000e-05, + 3.890870000000e-05, + 3.949570000000e-05, + 4.006100000000e-05, + 4.060510000000e-05,  \
+ 4.112870000000e-05, + 4.163230000000e-05, + 4.211650000000e-05, + 4.258190000000e-05, + 4.302910000000e-05,  \
+ 4.345860000000e-05, + 4.387110000000e-05, + 4.426700000000e-05, + 4.464700000000e-05, + 4.501150000000e-05 ]

.param id_pred_data_vd0.24=[ \
+ 3.516868396503e-10, + 5.052172546982e-10, + 7.323830075734e-10, + 1.065186232552e-09, + 1.549520618482e-09,  \
+ 2.252957287396e-09, + 3.276252016349e-09, + 4.768891841422e-09, + 6.949053812377e-09, + 1.012907347331e-08,  \
+ 1.474992075146e-08, + 2.143110521047e-08, + 3.104602569692e-08, + 4.483500674723e-08, + 6.456315077230e-08,  \
+ 9.272079296352e-08, + 1.327476411461e-07, + 1.892397176562e-07, + 2.680737270566e-07, + 3.763775475818e-07,  \
+ 5.222784602665e-07, + 7.144216397137e-07, + 9.613098882255e-07, + 1.270562606805e-06, + 1.648265133554e-06,  \
+ 2.098482800648e-06, + 2.623063555802e-06, + 3.221657389076e-06, + 3.891950327670e-06, + 4.630041948985e-06,  \
+ 5.430844612420e-06, + 6.288478762144e-06, + 7.196648803074e-06, + 8.148931665346e-06, + 9.138974128291e-06,  \
+ 1.016063906718e-05, + 1.120815955801e-05, + 1.227613189258e-05, + 1.335958979325e-05, + 1.445389701985e-05,  \
+ 1.555493508931e-05, + 1.665891031735e-05, + 1.776232849807e-05, + 1.886208134238e-05, + 1.995530154090e-05,  \
+ 2.103944483679e-05, + 2.211217302829e-05, + 2.317139238585e-05, + 2.421518904157e-05, + 2.524186740629e-05,  \
+ 2.624984190334e-05, + 2.723776444327e-05, + 2.820451743901e-05, + 2.914887503721e-05, + 3.007000079378e-05,  \
+ 3.096709144302e-05, + 3.183943452314e-05, + 3.268646774814e-05, + 3.350781393237e-05, + 3.430308192037e-05,  \
+ 3.507211105898e-05, + 3.581470227800e-05, + 3.653083811514e-05, + 3.722055698745e-05, + 3.788404050283e-05,  \
+ 3.852142137475e-05, + 3.913300693966e-05, + 3.971909754910e-05, + 4.028007388115e-05, + 4.081653314643e-05,  \
+ 4.132867092267e-05, + 4.181723808870e-05, + 4.228273755871e-05, + 4.272586433217e-05, + 4.314704448916e-05,  \
+ 4.354703938588e-05, + 4.392647766508e-05, + 4.428602987900e-05, + 4.462634562515e-05, + 4.494822816923e-05 ]

* Data table for Id-Vg at Vd = 0.25V
.param vg_data_vd0.25=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.25=[ \
+ 3.481190000000e-10, + 5.067510000000e-10, + 7.376500000000e-10, + 1.073700000000e-09, + 1.562800000000e-09,  \
+ 2.274500000000e-09, + 3.309900000000e-09, + 4.815900000000e-09, + 7.005400000000e-09, + 1.018670000000e-08,  \
+ 1.480520000000e-08, + 2.150190000000e-08, + 3.119450000000e-08, + 4.518810000000e-08, + 6.531850000000e-08,  \
+ 9.413120000000e-08, + 1.350850000000e-07, + 1.927530000000e-07, + 2.729620000000e-07, + 3.827910000000e-07,  \
+ 5.303500000000e-07, + 7.242790000000e-07, + 9.730300000000e-07, + 1.284100000000e-06, + 1.663200000000e-06,  \
+ 2.114000000000e-06, + 2.638000000000e-06, + 3.234500000000e-06, + 3.901100000000e-06, + 4.634200000000e-06,  \
+ 5.428900000000e-06, + 6.280100000000e-06, + 7.182300000000e-06, + 8.129900000000e-06, + 9.117300000000e-06,  \
+ 1.013930000000e-05, + 1.119050000000e-05, + 1.226610000000e-05, + 1.336120000000e-05, + 1.447130000000e-05,  \
+ 1.559200000000e-05, + 1.671920000000e-05, + 1.784880000000e-05, + 1.897720000000e-05, + 2.010070000000e-05,  \
+ 2.121620000000e-05, + 2.232070000000e-05, + 2.341130000000e-05, + 2.448570000000e-05, + 2.554160000000e-05,  \
+ 2.657720000000e-05, + 2.759100000000e-05, + 2.858160000000e-05, + 2.954800000000e-05, + 3.048940000000e-05,  \
+ 3.140530000000e-05, + 3.229530000000e-05, + 3.315930000000e-05, + 3.399700000000e-05, + 3.480870000000e-05,  \
+ 3.559450000000e-05, + 3.635460000000e-05, + 3.708950000000e-05, + 3.779940000000e-05, + 3.848480000000e-05,  \
+ 3.914620000000e-05, + 3.978400000000e-05, + 4.039890000000e-05, + 4.099120000000e-05, + 4.156170000000e-05,  \
+ 4.211090000000e-05, + 4.263930000000e-05, + 4.314740000000e-05, + 4.363600000000e-05, + 4.410560000000e-05,  \
+ 4.455670000000e-05, + 4.499000000000e-05, + 4.540590000000e-05, + 4.580510000000e-05, + 4.618800000000e-05 ]

.param id_pred_data_vd0.25=[ \
+ 3.551303140448e-10, + 5.100959099558e-10, + 7.395511425479e-10, + 1.075794342498e-09, + 1.565068519227e-09,  \
+ 2.275459154433e-09, + 3.308640028621e-09, + 4.815769116817e-09, + 7.017709968693e-09, + 1.023094320374e-08,  \
+ 1.490224121881e-08, + 2.165849366520e-08, + 3.138285009641e-08, + 4.532769892762e-08, + 6.527381657406e-08,  \
+ 9.373076181873e-08, + 1.341612403394e-07, + 1.911868565685e-07, + 2.707083410769e-07, + 3.798699879098e-07,  \
+ 5.268101403999e-07, + 7.201677476587e-07, + 9.684310953162e-07, + 1.279212028749e-06, + 1.658580572439e-06,  \
+ 2.110621380780e-06, + 2.637225179569e-06, + 3.238109002268e-06, + 3.911078692909e-06, + 4.652349616663e-06,  \
+ 5.456989583763e-06, + 6.319277417788e-06, + 7.233074484247e-06, + 8.192099812732e-06, + 9.190128366754e-06,  \
+ 1.022113792715e-05, + 1.127946597990e-05, + 1.235976014868e-05, + 1.345706550637e-05, + 1.456685731682e-05,  \
+ 1.568493462401e-05, + 1.680747845967e-05, + 1.793104456738e-05, + 1.905237877509e-05, + 2.016862708842e-05,  \
+ 2.127713923983e-05, + 2.237549233541e-05, + 2.346145993215e-05, + 2.453312845319e-05, + 2.558860796853e-05,  \
+ 2.662631959538e-05, + 2.764477721939e-05, + 2.864266207325e-05, + 2.961871905427e-05, + 3.057206413359e-05,  \
+ 3.150167322019e-05, + 3.240680962335e-05, + 3.328686943860e-05, + 3.414130333113e-05, + 3.496967838146e-05,  \
+ 3.577165625757e-05, + 3.654717875179e-05, + 3.729588206625e-05, + 3.801791535807e-05, + 3.871340595651e-05,  \
+ 3.938231020584e-05, + 4.002493005828e-05, + 4.064158565598e-05, + 4.123265171074e-05, + 4.179845564067e-05,  \
+ 4.233951040078e-05, + 4.285612521926e-05, + 4.334918412496e-05, + 4.381898907013e-05, + 4.426626765053e-05,  \
+ 4.469167834031e-05, + 4.509566861088e-05, + 4.547914431896e-05, + 4.584261841956e-05, + 4.618688035407e-05 ]

* Data table for Id-Vg at Vd = 0.26V
.param vg_data_vd0.26=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.26=[ \
+ 3.518670000000e-10, + 5.121430000000e-10, + 7.454050000000e-10, + 1.084900000000e-09, + 1.578800000000e-09,  \
+ 2.297600000000e-09, + 3.343100000000e-09, + 4.863500000000e-09, + 7.073700000000e-09, + 1.028470000000e-08,  \
+ 1.494560000000e-08, + 2.170290000000e-08, + 3.148170000000e-08, + 4.559740000000e-08, + 6.589980000000e-08,  \
+ 9.495300000000e-08, + 1.362400000000e-07, + 1.943620000000e-07, + 2.751780000000e-07, + 3.858070000000e-07,  \
+ 5.343890000000e-07, + 7.295950000000e-07, + 9.798980000000e-07, + 1.292800000000e-06, + 1.674000000000e-06,  \
+ 2.127300000000e-06, + 2.654000000000e-06, + 3.253600000000e-06, + 3.923600000000e-06, + 4.660400000000e-06,  \
+ 5.459300000000e-06, + 6.315100000000e-06, + 7.222500000000e-06, + 8.175900000000e-06, + 9.169800000000e-06,  \
+ 1.019910000000e-05, + 1.125860000000e-05, + 1.234360000000e-05, + 1.344920000000e-05, + 1.457110000000e-05,  \
+ 1.570500000000e-05, + 1.684690000000e-05, + 1.799280000000e-05, + 1.913910000000e-05, + 2.028240000000e-05,  \
+ 2.141920000000e-05, + 2.254670000000e-05, + 2.366190000000e-05, + 2.476240000000e-05, + 2.584580000000e-05,  \
+ 2.691020000000e-05, + 2.795370000000e-05, + 2.897490000000e-05, + 2.997260000000e-05, + 3.094590000000e-05,  \
+ 3.189390000000e-05, + 3.281620000000e-05, + 3.371240000000e-05, + 3.458230000000e-05, + 3.542580000000e-05,  \
+ 3.624320000000e-05, + 3.703440000000e-05, + 3.779990000000e-05, + 3.853980000000e-05, + 3.925470000000e-05,  \
+ 3.994490000000e-05, + 4.061090000000e-05, + 4.125310000000e-05, + 4.187230000000e-05, + 4.246870000000e-05,  \
+ 4.304310000000e-05, + 4.359600000000e-05, + 4.412790000000e-05, + 4.463940000000e-05, + 4.513120000000e-05,  \
+ 4.560370000000e-05, + 4.605750000000e-05, + 4.649330000000e-05, + 4.691150000000e-05, + 4.731280000000e-05 ]

.param id_pred_data_vd0.26=[ \
+ 3.585476271439e-10, + 5.149317283681e-10, + 7.466533702427e-10, + 1.086307985787e-09, + 1.580484338959e-09,  \
+ 2.297745282931e-09, + 3.340643726091e-09, + 4.861896485409e-09, + 7.085022986075e-09, + 1.033057422717e-08,  \
+ 1.505092207310e-08, + 2.188059127661e-08, + 3.171243747602e-08, + 4.581129530834e-08, + 6.597379979212e-08,  \
+ 9.472968486079e-08, + 1.355658207558e-07, + 1.931304416303e-07, + 2.733489782258e-07, + 3.833864002445e-07,  \
+ 5.313856081557e-07, + 7.259856283781e-07, + 9.756570034369e-07, + 1.287981449423e-06, + 1.669021075941e-06,  \
+ 2.122862297256e-06, + 2.651405138749e-06, + 3.254436305724e-06, + 3.929843423975e-06, + 4.673944204114e-06,  \
+ 5.481953230628e-06, + 6.348288661684e-06, + 7.266953180078e-06, + 8.231812316808e-06, + 9.236758560291e-06,  \
+ 1.027589911246e-05, + 1.134365142207e-05, + 1.243475169758e-05, + 1.354430693027e-05, + 1.466779584007e-05,  \
+ 1.580104712048e-05, + 1.694025268080e-05, + 1.808190048905e-05, + 1.922278592247e-05, + 2.035992758465e-05,  \
+ 2.149067324353e-05, + 2.261246714625e-05, + 2.372312243097e-05, + 2.482056384906e-05, + 2.590280695586e-05,  \
+ 2.696820025449e-05, + 2.801517170155e-05, + 2.904229302658e-05, + 3.004829675774e-05, + 3.103209703113e-05,  \
+ 3.199262311682e-05, + 3.292906912975e-05, + 3.384067269508e-05, + 3.472686628811e-05, + 3.558716183761e-05,  \
+ 3.642101451987e-05, + 3.722832596395e-05, + 3.800881240750e-05, + 3.876242466504e-05, + 3.948911733460e-05,  \
+ 4.018901527161e-05, + 4.086233035196e-05, + 4.150918364758e-05, + 4.212993837427e-05, + 4.272496153135e-05,  \
+ 4.329468443757e-05, + 4.383946652524e-05, + 4.435995477252e-05, + 4.485675453907e-05, + 4.533027065918e-05,  \
+ 4.578114254400e-05, + 4.621009284165e-05, + 4.661776096327e-05, + 4.700481280452e-05, + 4.737184615806e-05 ]

* Data table for Id-Vg at Vd = 0.27V
.param vg_data_vd0.27=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.27=[ \
+ 3.556230000000e-10, + 5.175460000000e-10, + 7.531760000000e-10, + 1.096000000000e-09, + 1.594900000000e-09,  \
+ 2.320600000000e-09, + 3.376200000000e-09, + 4.911100000000e-09, + 7.142000000000e-09, + 1.038270000000e-08,  \
+ 1.508600000000e-08, + 2.190370000000e-08, + 3.176860000000e-08, + 4.600610000000e-08, + 6.647990000000e-08,  \
+ 9.577260000000e-08, + 1.373900000000e-07, + 1.959630000000e-07, + 2.773840000000e-07, + 3.888040000000e-07,  \
+ 5.383990000000e-07, + 7.348650000000e-07, + 9.866960000000e-07, + 1.301400000000e-06, + 1.684700000000e-06,  \
+ 2.140300000000e-06, + 2.669700000000e-06, + 3.272200000000e-06, + 3.945500000000e-06, + 4.685800000000e-06,  \
+ 5.488600000000e-06, + 6.348800000000e-06, + 7.261000000000e-06, + 8.219700000000e-06, + 9.219700000000e-06,  \
+ 1.025570000000e-05, + 1.132270000000e-05, + 1.241610000000e-05, + 1.353120000000e-05, + 1.466370000000e-05,  \
+ 1.580950000000e-05, + 1.696450000000e-05, + 1.812510000000e-05, + 1.928760000000e-05, + 2.044860000000e-05,  \
+ 2.160470000000e-05, + 2.275310000000e-05, + 2.389070000000e-05, + 2.501510000000e-05, + 2.612380000000e-05,  \
+ 2.721480000000e-05, + 2.828600000000e-05, + 2.933590000000e-05, + 3.036320000000e-05, + 3.136660000000e-05,  \
+ 3.234520000000e-05, + 3.329840000000e-05, + 3.422570000000e-05, + 3.512670000000e-05, + 3.600120000000e-05,  \
+ 3.684920000000e-05, + 3.767080000000e-05, + 3.846610000000e-05, + 3.923550000000e-05, + 3.997930000000e-05,  \
+ 4.069780000000e-05, + 4.139140000000e-05, + 4.206070000000e-05, + 4.270620000000e-05, + 4.332820000000e-05,  \
+ 4.392750000000e-05, + 4.450460000000e-05, + 4.505990000000e-05, + 4.559410000000e-05, + 4.610770000000e-05,  \
+ 4.660140000000e-05, + 4.707570000000e-05, + 4.753110000000e-05, + 4.796820000000e-05, + 4.838770000000e-05 ]

.param id_pred_data_vd0.27=[ \
+ 3.619549160394e-10, + 5.197448271765e-10, + 7.537186474948e-10, + 1.096771313769e-09, + 1.595814160815e-09,  \
+ 2.319886283075e-09, + 3.372351358166e-09, + 4.907406641053e-09, + 7.151138241568e-09, + 1.042803059903e-08,  \
+ 1.519606648515e-08, + 2.209728720004e-08, + 3.203426643950e-08, + 4.628450071209e-08, + 6.666099352515e-08,  \
+ 9.571384197216e-08, + 1.369552995811e-07, + 1.950604286094e-07, + 2.759826952570e-07, + 3.869061231399e-07,  \
+ 5.359849114939e-07, + 7.318496068365e-07, + 9.829525379246e-07, + 1.296850309700e-06, + 1.679576357674e-06,  \
+ 2.135198319593e-06, + 2.665640186024e-06, + 3.270717170381e-06, + 3.948381026930e-06, + 4.695056104538e-06,  \
+ 5.506058278115e-06, + 6.375947086781e-06, + 7.298851105588e-06, + 8.268781530205e-06, + 9.279727455578e-06,  \
+ 1.032596675941e-05, + 1.140194381151e-05, + 1.250254990737e-05, + 1.362286886433e-05, + 1.475849036069e-05,  \
+ 1.590523981577e-05, + 1.705934046186e-05, + 1.821724734327e-05, + 1.937568857102e-05, + 2.053179989161e-05,  \
+ 2.168277795136e-05, + 2.282602566993e-05, + 2.395930154307e-05, + 2.508041317924e-05, + 2.618744321808e-05,  \
+ 2.727853716351e-05, + 2.835207233147e-05, + 2.940654587292e-05, + 3.044066514121e-05, + 3.145314534777e-05,  \
+ 3.244288047426e-05, + 3.340904149809e-05, + 3.435079546762e-05, + 3.526726621203e-05, + 3.615811583586e-05,  \
+ 3.702271176735e-05, + 3.786075933021e-05, + 3.867198349326e-05, + 3.945619959268e-05, + 4.021341941552e-05,  \
+ 4.094360760064e-05, + 4.164687808952e-05, + 4.232346269418e-05, + 4.297352250433e-05, + 4.359750542790e-05,  \
+ 4.419563541887e-05, + 4.476839967538e-05, + 4.531642291113e-05, + 4.584006266668e-05, + 4.633982185624e-05,  \
+ 4.681644699303e-05, + 4.727051564259e-05, + 4.770268395077e-05, + 4.811346661882e-05, + 4.850363766309e-05 ]

* Data table for Id-Vg at Vd = 0.28V
.param vg_data_vd0.28=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.28=[ \
+ 3.593920000000e-10, + 5.229650000000e-10, + 7.609670000000e-10, + 1.107200000000e-09, + 1.611000000000e-09,  \
+ 2.343800000000e-09, + 3.409400000000e-09, + 4.958800000000e-09, + 7.210400000000e-09, + 1.048070000000e-08,  \
+ 1.522640000000e-08, + 2.210450000000e-08, + 3.205530000000e-08, + 4.641440000000e-08, + 6.705930000000e-08,  \
+ 9.659080000000e-08, + 1.385380000000e-07, + 1.975600000000e-07, + 2.795820000000e-07, + 3.917870000000e-07,  \
+ 5.423850000000e-07, + 7.400970000000e-07, + 9.934340000000e-07, + 1.309900000000e-06, + 1.695200000000e-06,  \
+ 2.153200000000e-06, + 2.685100000000e-06, + 3.290500000000e-06, + 3.966800000000e-06, + 4.710600000000e-06,  \
+ 5.517100000000e-06, + 6.381400000000e-06, + 7.298100000000e-06, + 8.261800000000e-06, + 9.267300000000e-06,  \
+ 1.030940000000e-05, + 1.138330000000e-05, + 1.248430000000e-05, + 1.360800000000e-05, + 1.475010000000e-05,  \
+ 1.590660000000e-05, + 1.707360000000e-05, + 1.824740000000e-05, + 1.942440000000e-05, + 2.060130000000e-05,  \
+ 2.177490000000e-05, + 2.294220000000e-05, + 2.410030000000e-05, + 2.524650000000e-05, + 2.637850000000e-05,  \
+ 2.749400000000e-05, + 2.859100000000e-05, + 2.966770000000e-05, + 3.072260000000e-05, + 3.175450000000e-05,  \
+ 3.276220000000e-05, + 3.374490000000e-05, + 3.470190000000e-05, + 3.563280000000e-05, + 3.653720000000e-05,  \
+ 3.741490000000e-05, + 3.826610000000e-05, + 3.909060000000e-05, + 3.988880000000e-05, + 4.066080000000e-05,  \
+ 4.140710000000e-05, + 4.212790000000e-05, + 4.282370000000e-05, + 4.349510000000e-05, + 4.414240000000e-05,  \
+ 4.476620000000e-05, + 4.536700000000e-05, + 4.594540000000e-05, + 4.650200000000e-05, + 4.703730000000e-05,  \
+ 4.755190000000e-05, + 4.804630000000e-05, + 4.852110000000e-05, + 4.897690000000e-05, + 4.941430000000e-05 ]

.param id_pred_data_vd0.28=[ \
+ 3.653627578259e-10, + 5.245532097575e-10, + 7.607729202164e-10, + 1.107213698504e-09, + 1.611109290423e-09,  \
+ 2.341942426654e-09, + 3.403836110749e-09, + 4.952429222271e-09, + 7.216222570605e-09, + 1.052352047282e-08,  \
+ 1.533779297347e-08, + 2.230856949836e-08, + 3.234808559682e-08, + 4.674660942783e-08, + 6.733354211974e-08,  \
+ 9.668025427345e-08, + 1.383243943565e-07, + 1.969698155335e-07, + 2.785970218611e-07, + 3.904129289367e-07,  \
+ 5.405830506788e-07, + 7.377318434010e-07, + 9.902900001180e-07, + 1.305782298004e-06, + 1.690214030532e-06,  \
+ 2.147627710656e-06, + 2.679942954273e-06, + 3.286999963166e-06, + 3.966792537540e-06, + 4.715838222182e-06,  \
+ 5.529550107894e-06, + 6.402600993169e-06, + 7.329243744607e-06, + 8.303600843647e-06, + 9.319817181677e-06,  \
+ 1.037223832100e-05, + 1.145542832091e-05, + 1.256433679373e-05, + 1.369416189846e-05, + 1.484050924773e-05,  \
+ 1.599927578354e-05, + 1.716661616229e-05, + 1.833911490394e-05, + 1.951347367140e-05, + 2.068666100968e-05,  \
+ 2.185596938943e-05, + 2.301877480932e-05, + 2.417272829916e-05, + 2.531562960939e-05, + 2.644544758368e-05,  \
+ 2.756032423349e-05, + 2.865855843993e-05, + 2.973854891025e-05, + 3.079888178036e-05, + 3.183830209309e-05,  \
+ 3.285559971118e-05, + 3.384983341675e-05, + 3.482004976831e-05, + 3.576543997042e-05, + 3.668538469356e-05,  \
+ 3.757939091884e-05, + 3.844690450933e-05, + 3.928777063265e-05, + 4.010171629488e-05, + 4.088848072570e-05,  \
+ 4.164815763943e-05, + 4.238070629071e-05, + 4.308634262998e-05, + 4.376527038403e-05, + 4.441768920515e-05,  \
+ 4.504394950345e-05, + 4.564446688164e-05, + 4.621965286788e-05, + 4.677004937548e-05, + 4.729609237984e-05,  \
+ 4.779850714840e-05, + 4.827770520933e-05, + 4.873446479905e-05, + 4.916927486192e-05, + 4.958294623066e-05 ]

* Data table for Id-Vg at Vd = 0.29V
.param vg_data_vd0.29=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.29=[ \
+ 3.631750000000e-10, + 5.284040000000e-10, + 7.687830000000e-10, + 1.118500000000e-09, + 1.627100000000e-09,  \
+ 2.366900000000e-09, + 3.442700000000e-09, + 5.006500000000e-09, + 7.278900000000e-09, + 1.057890000000e-08,  \
+ 1.536700000000e-08, + 2.230550000000e-08, + 3.234210000000e-08, + 4.682260000000e-08, + 6.763840000000e-08,  \
+ 9.740810000000e-08, + 1.396850000000e-07, + 1.991540000000e-07, + 2.817720000000e-07, + 3.947590000000e-07,  \
+ 5.463510000000e-07, + 7.452960000000e-07, + 1.000100000000e-06, + 1.318300000000e-06, + 1.705700000000e-06,  \
+ 2.165900000000e-06, + 2.700300000000e-06, + 3.308400000000e-06, + 3.987800000000e-06, + 4.734800000000e-06,  \
+ 5.544900000000e-06, + 6.413000000000e-06, + 7.333900000000e-06, + 8.302300000000e-06, + 9.312900000000e-06,  \
+ 1.036070000000e-05, + 1.144090000000e-05, + 1.254900000000e-05, + 1.368050000000e-05, + 1.483130000000e-05,  \
+ 1.599740000000e-05, + 1.717520000000e-05, + 1.836090000000e-05, + 1.955110000000e-05, + 2.074250000000e-05,  \
+ 2.193190000000e-05, + 2.311630000000e-05, + 2.429300000000e-05, + 2.545920000000e-05, + 2.661250000000e-05,  \
+ 2.775060000000e-05, + 2.887140000000e-05, + 2.997300000000e-05, + 3.105380000000e-05, + 3.211240000000e-05,  \
+ 3.314760000000e-05, + 3.415820000000e-05, + 3.514360000000e-05, + 3.610320000000e-05, + 3.703630000000e-05,  \
+ 3.794280000000e-05, + 3.882260000000e-05, + 3.967550000000e-05, + 4.050170000000e-05, + 4.130140000000e-05,  \
+ 4.207480000000e-05, + 4.282230000000e-05, + 4.354420000000e-05, + 4.424100000000e-05, + 4.491310000000e-05,  \
+ 4.556110000000e-05, + 4.618540000000e-05, + 4.678660000000e-05, + 4.736520000000e-05, + 4.792180000000e-05,  \
+ 4.845700000000e-05, + 4.897130000000e-05, + 4.946530000000e-05, + 4.993950000000e-05, + 5.039460000000e-05 ]

.param id_pred_data_vd0.29=[ \
+ 3.687842653477e-10, + 5.293776383919e-10, + 7.678402291766e-10, + 1.117667665085e-09, + 1.626417058809e-09,  \
+ 2.363977733566e-09, + 3.435200834900e-09, + 4.997072604596e-09, + 7.280425489142e-09, + 1.061722979756e-08,  \
+ 1.547640827937e-08, + 2.251464884750e-08, + 3.265403670127e-08, + 4.719734292280e-08, + 6.799061921470e-08,  \
+ 9.762658891077e-08, + 1.396688992372e-07, + 1.988505937334e-07, + 2.811821605064e-07, + 3.938932138681e-07,  \
+ 5.451611991703e-07, + 7.436058103849e-07, + 9.976371893572e-07, + 1.314747846664e-06, + 1.700903885649e-06,  \
+ 2.160124513466e-06, + 2.694306513149e-06, + 3.303302974018e-06, + 3.985155790360e-06, + 4.736422451970e-06,  \
+ 5.552626535064e-06, + 6.428529632103e-06, + 7.358504299191e-06, + 8.336767477886e-06, + 9.357613125758e-06,  \
+ 1.041545547196e-05, + 1.150501258962e-05, + 1.262123623746e-05, + 1.375945797918e-05, + 1.491529634222e-05,  \
+ 1.608470323845e-05, + 1.726395552396e-05, + 1.844945349148e-05, + 1.963806796994e-05, + 2.082672886900e-05,  \
+ 2.201260242146e-05, + 2.319320512470e-05, + 2.436600916553e-05, + 2.552888130595e-05, + 2.667966509762e-05,  \
+ 2.781645518553e-05, + 2.893750446674e-05, + 3.004118399986e-05, + 3.112598722510e-05, + 3.219056583475e-05,  \
+ 3.323369601276e-05, + 3.425429742492e-05, + 3.525139945850e-05, + 3.622417920269e-05, + 3.717183906701e-05,  \
+ 3.809390007518e-05, + 3.898972077877e-05, + 3.985898889368e-05, + 4.070138369570e-05, + 4.151673638262e-05,  \
+ 4.230490347254e-05, + 4.306596092647e-05, + 4.379996360512e-05, + 4.450702967006e-05, + 4.518734902376e-05,  \
+ 4.584124661051e-05, + 4.646909801522e-05, + 4.707123662229e-05, + 4.764822369907e-05, + 4.820041373023e-05,  \
+ 4.872837220319e-05, + 4.923280386720e-05, + 4.971414760803e-05, + 5.017310395488e-05, + 5.061037765699e-05 ]

* Data table for Id-Vg at Vd = 0.30V
.param vg_data_vd0.30=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.30=[ \
+ 3.669740000000e-10, + 5.338630000000e-10, + 7.766290000000e-10, + 1.129700000000e-09, + 1.643300000000e-09,  \
+ 2.390200000000e-09, + 3.476100000000e-09, + 5.054400000000e-09, + 7.347500000000e-09, + 1.067720000000e-08,  \
+ 1.550780000000e-08, + 2.250670000000e-08, + 3.262920000000e-08, + 4.723110000000e-08, + 6.821750000000e-08,  \
+ 9.822520000000e-08, + 1.408300000000e-07, + 2.007450000000e-07, + 2.839580000000e-07, + 3.977210000000e-07,  \
+ 5.503000000000e-07, + 7.504670000000e-07, + 1.006800000000e-06, + 1.326700000000e-06, + 1.716000000000e-06,  \
+ 2.178400000000e-06, + 2.715300000000e-06, + 3.326100000000e-06, + 4.008300000000e-06, + 4.758500000000e-06,  \
+ 5.572000000000e-06, + 6.443800000000e-06, + 7.368700000000e-06, + 8.341500000000e-06, + 9.356800000000e-06,  \
+ 1.040990000000e-05, + 1.149600000000e-05, + 1.261050000000e-05, + 1.374910000000e-05, + 1.490790000000e-05,  \
+ 1.608290000000e-05, + 1.727040000000e-05, + 1.846690000000e-05, + 1.966900000000e-05, + 2.087350000000e-05,  \
+ 2.207730000000e-05, + 2.327730000000e-05, + 2.447090000000e-05, + 2.565530000000e-05, + 2.682810000000e-05,  \
+ 2.798700000000e-05, + 2.912970000000e-05, + 3.025440000000e-05, + 3.135940000000e-05, + 3.244300000000e-05,  \
+ 3.350400000000e-05, + 3.454110000000e-05, + 3.555350000000e-05, + 3.654030000000e-05, + 3.750110000000e-05,  \
+ 3.843520000000e-05, + 3.934260000000e-05, + 4.022310000000e-05, + 4.107660000000e-05, + 4.190320000000e-05,  \
+ 4.270320000000e-05, + 4.347670000000e-05, + 4.422420000000e-05, + 4.494600000000e-05, + 4.564250000000e-05,  \
+ 4.631420000000e-05, + 4.696160000000e-05, + 4.758520000000e-05, + 4.818550000000e-05, + 4.876310000000e-05,  \
+ 4.931860000000e-05, + 4.985250000000e-05, + 5.036540000000e-05, + 5.085790000000e-05, + 5.133050000000e-05 ]

.param id_pred_data_vd0.30=[ \
+ 3.722280150775e-10, + 5.342262965335e-10, + 7.749409780544e-10, + 1.128169158093e-09, + 1.641777114259e-09,  \
+ 2.386057484927e-09, + 3.466552112030e-09, + 5.041504813619e-09, + 7.343969699036e-09, + 1.070948876247e-08,  \
+ 1.561214304502e-08, + 2.271587931091e-08, + 3.295220736277e-08, + 4.763680436781e-08, + 6.863174775162e-08,  \
+ 9.855168627837e-08, + 1.409861965840e-07, + 2.006986960623e-07, + 2.837294005076e-07, + 3.973330422014e-07,  \
+ 5.497002234733e-07, + 7.494489636883e-07, + 1.004968362395e-06, + 1.323718606727e-06, + 1.711624599920e-06,  \
+ 2.172666108891e-06, + 2.708727151912e-06, + 3.319650295452e-06, + 4.003502817795e-06, + 4.756912312587e-06,  \
+ 5.575444993156e-06, + 6.453957394115e-06, + 7.386927063635e-06, + 8.368704948225e-06, + 9.393650179845e-06,  \
+ 1.045629323926e-05, + 1.155143363576e-05, + 1.267414372705e-05, + 1.381979927828e-05, + 1.498409255873e-05,  \
+ 1.616300723981e-05, + 1.735279984132e-05, + 1.855002265074e-05, + 1.975142440642e-05, + 2.095400050166e-05,  \
+ 2.215495915152e-05, + 2.335163517273e-05, + 2.454164714436e-05, + 2.572273588157e-05, + 2.689269458642e-05,  \
+ 2.804968753480e-05, + 2.919180042227e-05, + 3.031734813703e-05, + 3.142485729768e-05, + 3.251289599575e-05,  \
+ 3.358014364494e-05, + 3.462551321718e-05, + 3.564793296391e-05, + 3.664651012514e-05, + 3.762042179005e-05,  \
+ 3.856902185362e-05, + 3.949175588787e-05, + 4.038808256155e-05, + 4.125786654186e-05, + 4.210070183035e-05,  \
+ 4.291649238439e-05, + 4.370505484985e-05, + 4.446644161362e-05, + 4.520098445937e-05, + 4.590850876411e-05,  \
+ 4.658949910663e-05, + 4.724408208858e-05, + 4.787274228875e-05, + 4.847586824326e-05, + 4.905397508992e-05,  \
+ 4.960746009601e-05, + 5.013691261411e-05, + 5.064288707217e-05, + 5.112592043588e-05, + 5.158684652997e-05 ]

* Data table for Id-Vg at Vd = 0.31V
.param vg_data_vd0.31=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.31=[ \
+ 3.707900000000e-10, + 5.393470000000e-10, + 7.845060000000e-10, + 1.141100000000e-09, + 1.659600000000e-09,  \
+ 2.413500000000e-09, + 3.509500000000e-09, + 5.102400000000e-09, + 7.416400000000e-09, + 1.077580000000e-08,  \
+ 1.564880000000e-08, + 2.270830000000e-08, + 3.291670000000e-08, + 4.764000000000e-08, + 6.879700000000e-08,  \
+ 9.904250000000e-08, + 1.419740000000e-07, + 2.023340000000e-07, + 2.861400000000e-07, + 4.006750000000e-07,  \
+ 5.542360000000e-07, + 7.556150000000e-07, + 1.013400000000e-06, + 1.335000000000e-06, + 1.726300000000e-06,  \
+ 2.190800000000e-06, + 2.730100000000e-06, + 3.343500000000e-06, + 4.028500000000e-06, + 4.781700000000e-06,  \
+ 5.598500000000e-06, + 6.473800000000e-06, + 7.402500000000e-06, + 8.379400000000e-06, + 9.399300000000e-06,  \
+ 1.045730000000e-05, + 1.154880000000e-05, + 1.266920000000e-05, + 1.381450000000e-05, + 1.498050000000e-05,  \
+ 1.616360000000e-05, + 1.736000000000e-05, + 1.856630000000e-05, + 1.977930000000e-05, + 2.099570000000e-05,  \
+ 2.221250000000e-05, + 2.342680000000e-05, + 2.463580000000e-05, + 2.583690000000e-05, + 2.702750000000e-05,  \
+ 2.820540000000e-05, + 2.936840000000e-05, + 3.051450000000e-05, + 3.164190000000e-05, + 3.274880000000e-05,  \
+ 3.383400000000e-05, + 3.489600000000e-05, + 3.593390000000e-05, + 3.694670000000e-05, + 3.793380000000e-05,  \
+ 3.889450000000e-05, + 3.982850000000e-05, + 4.073550000000e-05, + 4.161550000000e-05, + 4.246830000000e-05,  \
+ 4.329410000000e-05, + 4.409320000000e-05, + 4.486570000000e-05, + 4.561190000000e-05, + 4.633240000000e-05,  \
+ 4.702740000000e-05, + 4.769750000000e-05, + 4.834310000000e-05, + 4.896490000000e-05, + 4.956320000000e-05,  \
+ 5.013870000000e-05, + 5.069190000000e-05, + 5.122340000000e-05, + 5.173380000000e-05, + 5.222360000000e-05 ]

.param id_pred_data_vd0.31=[ \
+ 3.757040478725e-10, + 5.391164148438e-10, + 7.820941472225e-10, + 1.138734941897e-09, + 1.657228776430e-09,  \
+ 2.408243142682e-09, + 3.497969913724e-09, + 5.085828647111e-09, + 7.407039124274e-09, + 1.080051323044e-08,  \
+ 1.574537680682e-08, + 2.291266660848e-08, + 3.324318576858e-08, + 4.806501635812e-08, + 6.925700247962e-08,  \
+ 9.945464711336e-08, + 1.422741601687e-07, + 2.025097461456e-07, + 2.862323503905e-07, + 4.007227460079e-07,  \
+ 5.541868415548e-07, + 7.552417423540e-07, + 1.012259122035e-06, + 1.332663218818e-06, + 1.722337697174e-06,  \
+ 2.185224689129e-06, + 2.723176421568e-06, + 3.336031622894e-06, + 4.021869835924e-06, + 4.777345802722e-06,  \
+ 5.598086863756e-06, + 6.479054409283e-06, + 7.414796218654e-06, + 8.399741655012e-06, + 9.428352786927e-06,  \
+ 1.049529186275e-05, + 1.159542469395e-05, + 1.272390185477e-05, + 1.387615924614e-05, + 1.504796997324e-05,  \
+ 1.623533269594e-05, + 1.743463853927e-05, + 1.864236095571e-05, + 1.985525195778e-05, + 2.107037820679e-05,  \
+ 2.228493380244e-05, + 2.349627073272e-05, + 2.470194398484e-05, + 2.589958974568e-05, + 2.708714644541e-05,  \
+ 2.826263822499e-05, + 2.942410952528e-05, + 3.056989575271e-05, + 3.169844960212e-05, + 3.280822376837e-05,  \
+ 3.389793033421e-05, + 3.496639641526e-05, + 3.601251453802e-05, + 3.703528775077e-05, + 3.803389729001e-05,  \
+ 3.900764844730e-05, + 3.995584876975e-05, + 4.087810579222e-05, + 4.177389622782e-05, + 4.264304865501e-05,  \
+ 4.348510294221e-05, + 4.430020795553e-05, + 4.508821482887e-05, + 4.584915965097e-05, + 4.658321835450e-05,  \
+ 4.729049469461e-05, + 4.797134955879e-05, + 4.862600850174e-05, + 4.925496774376e-05, + 4.985848441720e-05,  \
+ 5.043710887549e-05, + 5.099141402752e-05, + 5.152187804924e-05, + 5.202902422752e-05, + 5.251346156001e-05 ]

* Data table for Id-Vg at Vd = 0.32V
.param vg_data_vd0.32=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.32=[ \
+ 3.746240000000e-10, + 5.448560000000e-10, + 7.924190000000e-10, + 1.152400000000e-09, + 1.675900000000e-09,  \
+ 2.436900000000e-09, + 3.543100000000e-09, + 5.150600000000e-09, + 7.485400000000e-09, + 1.087470000000e-08,  \
+ 1.579020000000e-08, + 2.291030000000e-08, + 3.320470000000e-08, + 4.804960000000e-08, + 6.937720000000e-08,  \
+ 9.986030000000e-08, + 1.431190000000e-07, + 2.039230000000e-07, + 2.883200000000e-07, + 4.036250000000e-07,  \
+ 5.581610000000e-07, + 7.607440000000e-07, + 1.019900000000e-06, + 1.343200000000e-06, + 1.736400000000e-06,  \
+ 2.203100000000e-06, + 2.744800000000e-06, + 3.360600000000e-06, + 4.048500000000e-06, + 4.804500000000e-06,  \
+ 5.624400000000e-06, + 6.503200000000e-06, + 7.435500000000e-06, + 8.416300000000e-06, + 9.440400000000e-06,  \
+ 1.050300000000e-05, + 1.159950000000e-05, + 1.272550000000e-05, + 1.387690000000e-05, + 1.504970000000e-05,  \
+ 1.624010000000e-05, + 1.744470000000e-05, + 1.866010000000e-05, + 1.988290000000e-05, + 2.111020000000e-05,  \
+ 2.233890000000e-05, + 2.356610000000e-05, + 2.478920000000e-05, + 2.600550000000e-05, + 2.721250000000e-05,  \
+ 2.840790000000e-05, + 2.958960000000e-05, + 3.075540000000e-05, + 3.190350000000e-05, + 3.303220000000e-05,  \
+ 3.413990000000e-05, + 3.522540000000e-05, + 3.628730000000e-05, + 3.732470000000e-05, + 3.833680000000e-05,  \
+ 3.932290000000e-05, + 4.028240000000e-05, + 4.121500000000e-05, + 4.212050000000e-05, + 4.299870000000e-05,  \
+ 4.384970000000e-05, + 4.467360000000e-05, + 4.547050000000e-05, + 4.624070000000e-05, + 4.698460000000e-05,  \
+ 4.770250000000e-05, + 4.839490000000e-05, + 4.906230000000e-05, + 4.970510000000e-05, + 5.032380000000e-05,  \
+ 5.091900000000e-05, + 5.149120000000e-05, + 5.204110000000e-05, + 5.256910000000e-05, + 5.307580000000e-05 ]

.param id_pred_data_vd0.32=[ \
+ 3.792177238893e-10, + 5.440597306006e-10, + 7.893166298345e-10, + 1.149402137912e-09, + 1.672807314890e-09,  \
+ 2.430593895042e-09, + 3.529545722358e-09, + 5.130231102157e-09, + 7.469853926523e-09, + 1.089065335691e-08,  \
+ 1.587660335645e-08, + 2.310552190465e-08, + 3.352753310537e-08, + 4.848289336223e-08, + 6.986665539443e-08,  \
+ 1.003355737339e-07, + 1.435325793864e-07, + 2.042820597126e-07, + 2.886864422180e-07, + 4.040547719342e-07,  \
+ 5.586089537246e-07, + 7.609676686116e-07, + 1.019484407152e-06, + 1.341553579550e-06, + 1.733015960781e-06,  \
+ 2.197772701038e-06, + 2.737641043495e-06, + 3.352437051944e-06, + 4.040256899316e-06, + 4.797777510248e-06,  \
+ 5.620672018267e-06, + 6.503959302790e-06, + 7.442276109941e-06, + 8.430139860138e-06, + 9.462112793699e-06,  \
+ 1.053292304277e-05, + 1.163752167486e-05, + 1.277115428820e-05, + 1.392933889292e-05, + 1.510787289590e-05,  \
+ 1.630287035368e-05, + 1.751062110998e-05, + 1.872773165815e-05, + 1.995104830712e-05, + 2.117754891515e-05,  \
+ 2.240441506729e-05, + 2.362900413573e-05, + 2.484885742888e-05, + 2.606167690828e-05, + 2.726527396590e-05,  \
+ 2.845774870366e-05, + 2.963701495901e-05, + 3.080143127590e-05, + 3.194934688509e-05, + 3.307929029688e-05,  \
+ 3.418983658776e-05, + 3.527981461957e-05, + 3.634799504653e-05, + 3.739348612726e-05, + 3.841530531645e-05,  \
+ 3.941272851080e-05, + 4.038502462208e-05, + 4.133169073611e-05, + 4.225224256516e-05, + 4.314632620662e-05,  \
+ 4.401372279972e-05, + 4.485417157412e-05, + 4.566770978272e-05, + 4.645424894989e-05, + 4.721384029835e-05,  \
+ 4.794664680958e-05, + 4.865300375968e-05, + 4.933309741318e-05, + 4.998712334782e-05, + 5.061563104391e-05,  \
+ 5.121911410242e-05, + 5.179791245610e-05, + 5.235249176621e-05, + 5.288349930197e-05, + 5.339147057384e-05 ]

* Data table for Id-Vg at Vd = 0.33V
.param vg_data_vd0.33=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.33=[ \
+ 3.784790000000e-10, + 5.503920000000e-10, + 8.003700000000e-10, + 1.163800000000e-09, + 1.692300000000e-09,  \
+ 2.460400000000e-09, + 3.576800000000e-09, + 5.198900000000e-09, + 7.554600000000e-09, + 1.097380000000e-08,  \
+ 1.593200000000e-08, + 2.311290000000e-08, + 3.349340000000e-08, + 4.845990000000e-08, + 6.995830000000e-08,  \
+ 1.006790000000e-07, + 1.442650000000e-07, + 2.055120000000e-07, + 2.904990000000e-07, + 4.065700000000e-07,  \
+ 5.620780000000e-07, + 7.658560000000e-07, + 1.026500000000e-06, + 1.351400000000e-06, + 1.746500000000e-06,  \
+ 2.215300000000e-06, + 2.759200000000e-06, + 3.377600000000e-06, + 4.068100000000e-06, + 4.827000000000e-06,  \
+ 5.650000000000e-06, + 6.531900000000e-06, + 7.467700000000e-06, + 8.452200000000e-06, + 9.480400000000e-06,  \
+ 1.054740000000e-05, + 1.164860000000e-05, + 1.277980000000e-05, + 1.393680000000e-05, + 1.511580000000e-05,  \
+ 1.631310000000e-05, + 1.752520000000e-05, + 1.874880000000e-05, + 1.998070000000e-05, + 2.121790000000e-05,  \
+ 2.245750000000e-05, + 2.369660000000e-05, + 2.493250000000e-05, + 2.616270000000e-05, + 2.738480000000e-05,  \
+ 2.859630000000e-05, + 2.979510000000e-05, + 3.097910000000e-05, + 3.214640000000e-05, + 3.329530000000e-05,  \
+ 3.442410000000e-05, + 3.553150000000e-05, + 3.661600000000e-05, + 3.767660000000e-05, + 3.871240000000e-05,  \
+ 3.972260000000e-05, + 4.070650000000e-05, + 4.166370000000e-05, + 4.259370000000e-05, + 4.349650000000e-05,  \
+ 4.437190000000e-05, + 4.521990000000e-05, + 4.604060000000e-05, + 4.683420000000e-05, + 4.760110000000e-05,  \
+ 4.834150000000e-05, + 4.905580000000e-05, + 4.974440000000e-05, + 5.040790000000e-05, + 5.104660000000e-05,  \
+ 5.166120000000e-05, + 5.225220000000e-05, + 5.282010000000e-05, + 5.336550000000e-05, + 5.388890000000e-05 ]

.param id_pred_data_vd0.33=[ \
+ 3.827742756091e-10, + 5.490627885685e-10, + 7.966236270640e-10, + 1.160186480220e-09, + 1.688557293988e-09,  \
+ 2.453155838467e-09, + 3.561350681025e-09, + 5.174801387398e-09, + 7.532623591544e-09, + 1.098015694367e-08,  \
+ 1.600616844399e-08, + 2.329505804255e-08, + 3.380591444113e-08, + 4.889109234796e-08, + 7.046167382896e-08,  \
+ 1.011953938246e-07, + 1.447614704375e-07, + 2.060145590121e-07, + 2.910900866482e-07, + 4.073237789726e-07,  \
+ 5.629576889987e-07, + 7.666131068618e-07, + 1.026632498906e-06, + 1.350373781861e-06, + 1.743643033478e-06,  \
+ 2.210284210378e-06, + 2.752097061602e-06, + 3.368863990545e-06, + 4.058671947860e-06, + 4.818220368179e-06,  \
+ 5.643238055200e-06, + 6.528770409204e-06, + 7.469533884432e-06, + 8.460127883154e-06, + 9.495192625764e-06,  \
+ 1.056954421074e-05, + 1.167821723357e-05, + 1.281649900193e-05, + 1.398002197675e-05, + 1.516460950370e-05,  \
+ 1.636643428355e-05, + 1.758186230290e-05, + 1.880751166027e-05, + 2.004018653679e-05, + 2.127693602233e-05,  \
+ 2.251494726806e-05, + 2.375158030191e-05, + 2.498440764612e-05, + 2.621104264108e-05, + 2.742935554124e-05,  \
+ 2.863728142984e-05, + 2.983289225085e-05, + 3.101446643996e-05, + 3.218020079657e-05, + 3.332876753120e-05,  \
+ 3.445859634667e-05, + 3.556850351742e-05, + 3.665727410407e-05, + 3.772396448767e-05, + 3.876741735439e-05,  \
+ 3.978699642175e-05, + 4.078198136995e-05, + 4.175164227490e-05, + 4.269564058632e-05, + 4.361345287180e-05,  \
+ 4.450483422261e-05, + 4.536950131296e-05, + 4.620749736205e-05, + 4.701849102275e-05, + 4.780275601661e-05,  \
+ 4.856031155214e-05, + 4.929116723360e-05, + 4.999591372325e-05, + 5.067447898909e-05, + 5.132743928698e-05,  \
+ 5.195511155762e-05, + 5.255786556518e-05, + 5.313629197190e-05, + 5.369086138671e-05, + 5.422209724202e-05 ]

* Data table for Id-Vg at Vd = 0.34V
.param vg_data_vd0.34=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.34=[ \
+ 3.823550000000e-10, + 5.559580000000e-10, + 8.083600000000e-10, + 1.175300000000e-09, + 1.708700000000e-09,  \
+ 2.484000000000e-09, + 3.610700000000e-09, + 5.247400000000e-09, + 7.624200000000e-09, + 1.107330000000e-08,  \
+ 1.607430000000e-08, + 2.331600000000e-08, + 3.378280000000e-08, + 4.887120000000e-08, + 7.054050000000e-08,  \
+ 1.014990000000e-07, + 1.454120000000e-07, + 2.071020000000e-07, + 2.926780000000e-07, + 4.095130000000e-07,  \
+ 5.659880000000e-07, + 7.709540000000e-07, + 1.033000000000e-06, + 1.359600000000e-06, + 1.756500000000e-06,  \
+ 2.227400000000e-06, + 2.773600000000e-06, + 3.394400000000e-06, + 4.087500000000e-06, + 4.849200000000e-06,  \
+ 5.675000000000e-06, + 6.560100000000e-06, + 7.499300000000e-06, + 8.487300000000e-06, + 9.519300000000e-06,  \
+ 1.059040000000e-05, + 1.169610000000e-05, + 1.283210000000e-05, + 1.399440000000e-05, + 1.517920000000e-05,  \
+ 1.638280000000e-05, + 1.760190000000e-05, + 1.883310000000e-05, + 2.007340000000e-05, + 2.131970000000e-05,  \
+ 2.256920000000e-05, + 2.381920000000e-05, + 2.506690000000e-05, + 2.630990000000e-05, + 2.754570000000e-05,  \
+ 2.877200000000e-05, + 2.998660000000e-05, + 3.118740000000e-05, + 3.237250000000e-05, + 3.354010000000e-05,  \
+ 3.468860000000e-05, + 3.581640000000e-05, + 3.692210000000e-05, + 3.800460000000e-05, + 3.906280000000e-05,  \
+ 4.009580000000e-05, + 4.110290000000e-05, + 4.208360000000e-05, + 4.303720000000e-05, + 4.396360000000e-05,  \
+ 4.486250000000e-05, + 4.573390000000e-05, + 4.657780000000e-05, + 4.739420000000e-05, + 4.818350000000e-05,  \
+ 4.894590000000e-05, + 4.968160000000e-05, + 5.039120000000e-05, + 5.107500000000e-05, + 5.173340000000e-05,  \
+ 5.236710000000e-05, + 5.297650000000e-05, + 5.356220000000e-05, + 5.412470000000e-05, + 5.466460000000e-05 ]

.param id_pred_data_vd0.34=[ \
+ 3.863791997460e-10, + 5.541333836234e-10, + 8.040263832498e-10, + 1.171101695618e-09, + 1.704495575794e-09,  \
+ 2.475980522831e-09, + 3.593485633502e-09, + 5.219682002178e-09, + 7.595519697645e-09, + 1.106938988471e-08,  \
+ 1.613452361937e-08, + 2.348186171730e-08, + 3.407934642041e-08, + 4.929081541150e-08, + 7.104344888376e-08,  \
+ 1.020351976422e-07, + 1.459612951749e-07, + 2.077076146634e-07, + 2.934411520528e-07, + 4.105279163014e-07,  \
+ 5.672286101799e-07, + 7.721720339759e-07, + 1.033684466165e-06, + 1.359103853247e-06, + 1.754186014296e-06,  \
+ 2.222743423772e-06, + 2.766517809505e-06, + 3.385282816453e-06, + 4.077103603777e-06, + 4.838707609451e-06,  \
+ 5.665817589033e-06, + 6.553554849233e-06, + 7.496681682824e-06, + 8.489879983244e-06, + 9.527830407023e-06,  \
+ 1.060546099325e-05, + 1.171786738269e-05, + 1.286041857384e-05, + 1.402879774105e-05, + 1.521888225398e-05,  \
+ 1.642690447625e-05, + 1.764929715137e-05, + 1.888261795102e-05, + 2.012384262343e-05, + 2.136987022823e-05,  \
+ 2.261805624585e-05, + 2.386567823123e-05, + 2.511024751584e-05, + 2.634954260429e-05, + 2.758126283879e-05,  \
+ 2.880337473471e-05, + 3.001399076311e-05, + 3.121125060716e-05, + 3.239346464397e-05, + 3.355917579029e-05,  \
+ 3.470687501249e-05, + 3.583523634006e-05, + 3.694316386827e-05, + 3.802941326285e-05, + 3.909309642040e-05,  \
+ 4.013344645500e-05, + 4.114960989682e-05, + 4.214095592033e-05, + 4.310694523156e-05, + 4.404712264659e-05,  \
+ 4.496117646340e-05, + 4.584891867125e-05, + 4.671002272516e-05, + 4.754452325869e-05, + 4.835236584768e-05,  \
+ 4.913352575386e-05, + 4.988828004571e-05, + 5.061676725745e-05, + 5.131907644682e-05, + 5.199581122724e-05,  \
+ 5.264706560411e-05, + 5.327339371433e-05, + 5.387510231230e-05, + 5.445280490676e-05, + 5.500689730980e-05 ]

* Data table for Id-Vg at Vd = 0.35V
.param vg_data_vd0.35=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.35=[ \
+ 3.862530000000e-10, + 5.615540000000e-10, + 8.163930000000e-10, + 1.186800000000e-09, + 1.725300000000e-09,  \
+ 2.507800000000e-09, + 3.644700000000e-09, + 5.296200000000e-09, + 7.693900000000e-09, + 1.117320000000e-08,  \
+ 1.621710000000e-08, + 2.351970000000e-08, + 3.407300000000e-08, + 4.928350000000e-08, + 7.112400000000e-08,  \
+ 1.023210000000e-07, + 1.465610000000e-07, + 2.086930000000e-07, + 2.948570000000e-07, + 4.124550000000e-07,  \
+ 5.698930000000e-07, + 7.760420000000e-07, + 1.039500000000e-06, + 1.367700000000e-06, + 1.766500000000e-06,  \
+ 2.239400000000e-06, + 2.787800000000e-06, + 3.411000000000e-06, + 4.106600000000e-06, + 4.871000000000e-06,  \
+ 5.699800000000e-06, + 6.587900000000e-06, + 7.530200000000e-06, + 8.521700000000e-06, + 9.557300000000e-06,  \
+ 1.063230000000e-05, + 1.174220000000e-05, + 1.288280000000e-05, + 1.405000000000e-05, + 1.524020000000e-05,  \
+ 1.644970000000e-05, + 1.767520000000e-05, + 1.891350000000e-05, + 2.016150000000e-05, + 2.141620000000e-05,  \
+ 2.267490000000e-05, + 2.393480000000e-05, + 2.519340000000e-05, + 2.644810000000e-05, + 2.769660000000e-05,  \
+ 2.893650000000e-05, + 3.016560000000e-05, + 3.138200000000e-05, + 3.258350000000e-05, + 3.376850000000e-05,  \
+ 3.493520000000e-05, + 3.608200000000e-05, + 3.720760000000e-05, + 3.831060000000e-05, + 3.938990000000e-05,  \
+ 4.044460000000e-05, + 4.147380000000e-05, + 4.247670000000e-05, + 4.345300000000e-05, + 4.440200000000e-05,  \
+ 4.532360000000e-05, + 4.621760000000e-05, + 4.708390000000e-05, + 4.792260000000e-05, + 4.873370000000e-05,  \
+ 4.951750000000e-05, + 5.027420000000e-05, + 5.100430000000e-05, + 5.170800000000e-05, + 5.238590000000e-05,  \
+ 5.303830000000e-05, + 5.366590000000e-05, + 5.426900000000e-05, + 5.484830000000e-05, + 5.540440000000e-05 ]

.param id_pred_data_vd0.35=[ \
+ 3.900331280171e-10, + 5.592744933836e-10, + 8.115293437250e-10, + 1.182167608249e-09, + 1.720644315917e-09,  \
+ 2.499104811982e-09, + 3.625995015355e-09, + 5.264995195375e-09, + 7.658769707319e-09, + 1.115860897016e-08,  \
+ 1.626217951411e-08, + 2.366656737252e-08, + 3.434832578364e-08, + 4.968307578679e-08, + 7.161284472090e-08,  \
+ 1.028563261229e-07, + 1.471347971460e-07, + 2.093631621847e-07, + 2.957414210414e-07, + 4.136662994370e-07,  \
+ 5.714188546335e-07, + 7.776359893796e-07, + 1.040636561811e-06, + 1.367729191770e-06, + 1.764635339896e-06,  \
+ 2.235124588879e-06, + 2.780893601084e-06, + 3.401683261472e-06, + 4.095558324479e-06, + 4.859228602072e-06,  \
+ 5.688446708518e-06, + 6.578374450328e-06, + 7.523817112087e-06, + 8.519505809090e-06, + 9.560229591443e-06,  \
+ 1.064093603418e-05, + 1.175681718451e-05, + 1.290331401833e-05, + 1.407613999618e-05, + 1.527128933958e-05,  \
+ 1.648494981055e-05, + 1.771365423338e-05, + 1.895403984236e-05, + 2.020300235017e-05, + 2.145757498511e-05,  \
+ 2.271493358421e-05, + 2.397263087914e-05, + 2.522799804865e-05, + 2.647880937729e-05, + 2.772278567136e-05,  \
+ 2.895796351368e-05, + 3.018232855538e-05, + 3.139402688248e-05, + 3.259136756242e-05, + 3.377289649507e-05,  \
+ 3.493703225104e-05, + 3.608251172409e-05, + 3.720805143530e-05, + 3.831257672573e-05, + 3.939510970667e-05,  \
+ 4.045468522236e-05, + 4.149061314820e-05, + 4.250221099937e-05, + 4.348888032837e-05, + 4.445015001693e-05,  \
+ 4.538567372947e-05, + 4.629508475773e-05, + 4.717824558611e-05, + 4.803494230146e-05, + 4.886519018328e-05,  \
+ 4.966908090864e-05, + 5.044654317317e-05, + 5.119787747390e-05, + 5.192315002205e-05, + 5.262285485514e-05,  \
+ 5.329695632099e-05, + 5.394613690441e-05, + 5.457064107759e-05, + 5.517100362340e-05, + 5.574755050475e-05 ]

* Data table for Id-Vg at Vd = 0.36V
.param vg_data_vd0.36=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.36=[ \
+ 3.901740000000e-10, + 5.671820000000e-10, + 8.244700000000e-10, + 1.198400000000e-09, + 1.741900000000e-09,  \
+ 2.531600000000e-09, + 3.678900000000e-09, + 5.345100000000e-09, + 7.764000000000e-09, + 1.127340000000e-08,  \
+ 1.636030000000e-08, + 2.372420000000e-08, + 3.436420000000e-08, + 4.969700000000e-08, + 7.170900000000e-08,  \
+ 1.031440000000e-07, + 1.477110000000e-07, + 2.102860000000e-07, + 2.970370000000e-07, + 4.153970000000e-07,  \
+ 5.737950000000e-07, + 7.811210000000e-07, + 1.046000000000e-06, + 1.375800000000e-06, + 1.776400000000e-06,  \
+ 2.251400000000e-06, + 2.802000000000e-06, + 3.427500000000e-06, + 4.125600000000e-06, + 4.892600000000e-06,  \
+ 5.724100000000e-06, + 6.615200000000e-06, + 7.560600000000e-06, + 8.555300000000e-06, + 9.594400000000e-06,  \
+ 1.067320000000e-05, + 1.178710000000e-05, + 1.293200000000e-05, + 1.410390000000e-05, + 1.529910000000e-05,  \
+ 1.651410000000e-05, + 1.774560000000e-05, + 1.899040000000e-05, + 2.024550000000e-05, + 2.150800000000e-05,  \
+ 2.277520000000e-05, + 2.404430000000e-05, + 2.531290000000e-05, + 2.657840000000e-05, + 2.783850000000e-05,  \
+ 2.909090000000e-05, + 3.033350000000e-05, + 3.156420000000e-05, + 3.278100000000e-05, + 3.398210000000e-05,  \
+ 3.516570000000e-05, + 3.633030000000e-05, + 3.747440000000e-05, + 3.859660000000e-05, + 3.969580000000e-05,  \
+ 4.077090000000e-05, + 4.182090000000e-05, + 4.284510000000e-05, + 4.384290000000e-05, + 4.481360000000e-05,  \
+ 4.575700000000e-05, + 4.667280000000e-05, + 4.756080000000e-05, + 4.842090000000e-05, + 4.925320000000e-05,  \
+ 5.005790000000e-05, + 5.083520000000e-05, + 5.158530000000e-05, + 5.230860000000e-05, + 5.300540000000e-05,  \
+ 5.367630000000e-05, + 5.432170000000e-05, + 5.494210000000e-05, + 5.553800000000e-05, + 5.611000000000e-05 ]

.param id_pred_data_vd0.36=[ \
+ 3.937402404119e-10, + 5.644933320781e-10, + 8.191473899188e-10, + 1.193396901300e-09, + 1.737031478655e-09,  \
+ 2.522554805040e-09, + 3.658965290754e-09, + 5.310821862281e-09, + 7.722529815624e-09, + 1.124811475961e-08,  \
+ 1.638946386606e-08, + 2.384980405168e-08, + 3.461413683681e-08, + 5.006908168070e-08, + 7.217198742637e-08,  \
+ 1.036613866745e-07, + 1.482831726207e-07, + 2.109833485520e-07, + 2.979933765346e-07, + 4.167399174548e-07,  \
+ 5.755284837505e-07, + 7.830046524759e-07, + 1.047481200658e-06, + 1.376246127620e-06, + 1.774978827598e-06,  \
+ 2.247411212011e-06, + 2.795201980916e-06, + 3.418057603994e-06, + 4.114017174288e-06, + 4.879779335170e-06,  \
+ 5.711142657674e-06, + 6.603247602470e-06, + 7.550990703749e-06, + 8.549126068829e-06, + 9.592489659553e-06,  \
+ 1.067614990461e-05, + 1.179530750960e-05, + 1.294547095313e-05, + 1.412243946106e-05, + 1.532223555841e-05,  \
+ 1.654114370467e-05, + 1.777566445526e-05, + 1.902249612613e-05, + 2.027856098721e-05, + 2.154092668206e-05,  \
+ 2.280684420839e-05, + 2.407364838291e-05, + 2.533892024076e-05, + 2.660033118445e-05, + 2.785562071949e-05,  \
+ 2.910271170549e-05, + 3.033970511751e-05, + 3.156473336276e-05, + 3.277605457697e-05, + 3.397208667593e-05,  \
+ 3.515143616823e-05, + 3.631267027231e-05, + 3.745453432202e-05, + 3.857597534079e-05, + 3.967590106186e-05,  \
+ 4.075344448211e-05, + 4.180778574664e-05, + 4.283822810976e-05, + 4.384423722513e-05, + 4.482528136577e-05,  \
+ 4.578079737257e-05, + 4.671068571042e-05, + 4.761457967106e-05, + 4.849242162891e-05, + 4.934403346851e-05,  \
+ 5.016938899644e-05, + 5.096858250909e-05, + 5.174175021239e-05, + 5.248909641523e-05, + 5.321073636878e-05,  \
+ 5.390712060034e-05, + 5.457830673549e-05, + 5.522497580387e-05, + 5.584729020484e-05, + 5.644592049066e-05 ]

* Data table for Id-Vg at Vd = 0.37V
.param vg_data_vd0.37=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.37=[ \
+ 3.941190000000e-10, + 5.728430000000e-10, + 8.325920000000e-10, + 1.210100000000e-09, + 1.758600000000e-09,  \
+ 2.555500000000e-09, + 3.713200000000e-09, + 5.394300000000e-09, + 7.834400000000e-09, + 1.137410000000e-08,  \
+ 1.650420000000e-08, + 2.392940000000e-08, + 3.465640000000e-08, + 5.011180000000e-08, + 7.229560000000e-08,  \
+ 1.039690000000e-07, + 1.488640000000e-07, + 2.118820000000e-07, + 2.992200000000e-07, + 4.183390000000e-07,  \
+ 5.776950000000e-07, + 7.861930000000e-07, + 1.052400000000e-06, + 1.383900000000e-06, + 1.786300000000e-06,  \
+ 2.263300000000e-06, + 2.816000000000e-06, + 3.443800000000e-06, + 4.144400000000e-06, + 4.914000000000e-06,  \
+ 5.748200000000e-06, + 6.642100000000e-06, + 7.590500000000e-06, + 8.588400000000e-06, + 9.630800000000e-06,  \
+ 1.071310000000e-05, + 1.183090000000e-05, + 1.297980000000e-05, + 1.415610000000e-05, + 1.535610000000e-05,  \
+ 1.657630000000e-05, + 1.781340000000e-05, + 1.906430000000e-05, + 2.032600000000e-05, + 2.159570000000e-05,  \
+ 2.287070000000e-05, + 2.414830000000e-05, + 2.542610000000e-05, + 2.670160000000e-05, + 2.797240000000e-05,  \
+ 2.923640000000e-05, + 3.049140000000e-05, + 3.173530000000e-05, + 3.296620000000e-05, + 3.418220000000e-05,  \
+ 3.538160000000e-05, + 3.656280000000e-05, + 3.772410000000e-05, + 3.886440000000e-05, + 3.998220000000e-05,  \
+ 4.107650000000e-05, + 4.214630000000e-05, + 4.319060000000e-05, + 4.420880000000e-05, + 4.520030000000e-05,  \
+ 4.616450000000e-05, + 4.710120000000e-05, + 4.801010000000e-05, + 4.889100000000e-05, + 4.974390000000e-05,  \
+ 5.056890000000e-05, + 5.136610000000e-05, + 5.213580000000e-05, + 5.287820000000e-05, + 5.359370000000e-05,  \
+ 5.428270000000e-05, + 5.494560000000e-05, + 5.558290000000e-05, + 5.619510000000e-05, + 5.678280000000e-05 ]

.param id_pred_data_vd0.37=[ \
+ 3.975002771384e-10, + 5.697905169910e-10, + 8.268767848207e-10, + 1.204793333986e-09, + 1.753666230009e-09,  \
+ 2.546367223744e-09, + 3.692413317324e-09, + 5.357264916128e-09, + 7.786928168940e-09, + 1.133812858711e-08,  \
+ 1.651684080173e-08, + 2.403232059578e-08, + 3.487743128971e-08, + 5.045022945183e-08, + 7.272249746393e-08,  \
+ 1.044521857807e-07, + 1.494099598176e-07, + 2.125711858980e-07, + 3.001999806429e-07, + 4.197533257866e-07,  \
+ 5.795607603432e-07, + 7.882799445724e-07, + 1.054219721937e-06, + 1.384645240705e-06, + 1.785210256458e-06,  \
+ 2.259598577439e-06, + 2.809432617141e-06, + 3.434388145251e-06, + 4.132466610827e-06, + 4.900373214696e-06,  \
+ 5.733894140576e-06, + 6.628219271079e-06, + 7.578230579384e-06, + 8.578788165323e-06, + 9.624771646486e-06,  \
+ 1.071124101145e-05, + 1.183351199870e-05, + 1.298716753809e-05, + 1.416802140739e-05, + 1.537217274745e-05,  \
+ 1.659592395299e-05, + 1.783584259101e-05, + 1.908866179292e-05, + 2.035126948613e-05, + 2.162084165320e-05,  \
+ 2.289455696882e-05, + 2.416987408651e-05, + 2.544425435190e-05, + 2.671539332368e-05, + 2.798110232106e-05,  \
+ 2.923921958427e-05, + 3.048786064028e-05, + 3.172510332661e-05, + 3.294927046227e-05, + 3.415875486098e-05,  \
+ 3.535213778378e-05, + 3.652787396277e-05, + 3.768491078517e-05, + 3.882195065671e-05, + 3.993799211457e-05,  \
+ 4.103220060642e-05, + 4.210367158521e-05, + 4.315165126172e-05, + 4.417563621246e-05, + 4.517503955867e-05,  \
+ 4.614940902684e-05, + 4.709846194601e-05, + 4.802189680049e-05, + 4.891951975878e-05, + 4.979130928405e-05,  \
+ 5.063708769740e-05, + 5.145687653567e-05, + 5.225085886195e-05, + 5.301920697093e-05, + 5.376202854677e-05,  \
+ 5.447954972624e-05, + 5.517212048289e-05, + 5.584015001659e-05, + 5.648377293255e-05, + 5.710366225685e-05 ]

* Data table for Id-Vg at Vd = 0.38V
.param vg_data_vd0.38=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.38=[ \
+ 3.980880000000e-10, + 5.785380000000e-10, + 8.407630000000e-10, + 1.221800000000e-09, + 1.775400000000e-09,  \
+ 2.579600000000e-09, + 3.747700000000e-09, + 5.443700000000e-09, + 7.905100000000e-09, + 1.147530000000e-08,  \
+ 1.664860000000e-08, + 2.413540000000e-08, + 3.494960000000e-08, + 5.052790000000e-08, + 7.288400000000e-08,  \
+ 1.047960000000e-07, + 1.500190000000e-07, + 2.134800000000e-07, + 3.014050000000e-07, + 4.212830000000e-07,  \
+ 5.815940000000e-07, + 7.912600000000e-07, + 1.058900000000e-06, + 1.392000000000e-06, + 1.796200000000e-06,  \
+ 2.275100000000e-06, + 2.830000000000e-06, + 3.460100000000e-06, + 4.163000000000e-06, + 4.935100000000e-06,  \
+ 5.772000000000e-06, + 6.668600000000e-06, + 7.619900000000e-06, + 8.620900000000e-06, + 9.666500000000e-06,  \
+ 1.075220000000e-05, + 1.187360000000e-05, + 1.302650000000e-05, + 1.420690000000e-05, + 1.541140000000e-05,  \
+ 1.663640000000e-05, + 1.787880000000e-05, + 1.913530000000e-05, + 2.040320000000e-05, + 2.167970000000e-05,  \
+ 2.296190000000e-05, + 2.424740000000e-05, + 2.553370000000e-05, + 2.681840000000e-05, + 2.809930000000e-05,  \
+ 2.937390000000e-05, + 3.064040000000e-05, + 3.189660000000e-05, + 3.314050000000e-05, + 3.437040000000e-05,  \
+ 3.558440000000e-05, + 3.678090000000e-05, + 3.795840000000e-05, + 3.911550000000e-05, + 4.025080000000e-05,  \
+ 4.136320000000e-05, + 4.245150000000e-05, + 4.351490000000e-05, + 4.455250000000e-05, + 4.556370000000e-05,  \
+ 4.654790000000e-05, + 4.750460000000e-05, + 4.843360000000e-05, + 4.933450000000e-05, + 5.020730000000e-05,  \
+ 5.105200000000e-05, + 5.186870000000e-05, + 5.265740000000e-05, + 5.341850000000e-05, + 5.415220000000e-05,  \
+ 5.485900000000e-05, + 5.553910000000e-05, + 5.619300000000e-05, + 5.682130000000e-05, + 5.742430000000e-05 ]

.param id_pred_data_vd0.38=[ \
+ 4.013137333558e-10, + 5.751690634881e-10, + 8.347267366204e-10, + 1.216365537182e-09, + 1.770564566073e-09,  \
+ 2.570560653226e-09, + 3.726386825775e-09, + 5.404401353104e-09, + 7.852147305698e-09, + 1.142892536166e-08,  \
+ 1.664472904395e-08, + 2.421456457569e-08, + 3.513930323606e-08, + 5.082767017939e-08, + 7.326600950819e-08,  \
+ 1.052311301919e-07, + 1.505180023287e-07, + 2.141308891623e-07, + 3.023663145996e-07, + 4.227106660437e-07,  \
+ 5.835192973791e-07, + 7.934643554108e-07, + 1.060851577677e-06, + 1.392931862938e-06, + 1.795325661078e-06,  \
+ 2.271680432386e-06, + 2.823579061442e-06, + 3.450661079114e-06, + 4.150895347266e-06, + 4.920991505060e-06,  \
+ 5.756712744187e-06, + 6.653283453488e-06, + 7.605618011439e-06, + 8.608576536062e-06, + 9.657104856160e-06,  \
+ 1.074633266398e-05, + 1.187162466522e-05, + 1.302860961005e-05, + 1.421316301276e-05, + 1.542138779769e-05,  \
+ 1.664970761340e-05, + 1.789465117326e-05, + 1.915302505950e-05, + 2.042176027317e-05, + 2.169804771256e-05,  \
+ 2.297902712598e-05, + 2.426217281027e-05, + 2.554497841629e-05, + 2.682516293135e-05, + 2.810044257785e-05,  \
+ 2.936879624031e-05, + 3.062817238970e-05, + 3.187676004018e-05, + 3.311284497613e-05, + 3.433475169004e-05,  \
+ 3.554102586349e-05, + 3.673025741591e-05, + 3.790122704231e-05, + 3.905272373231e-05, + 4.018371619168e-05,  \
+ 4.129331689910e-05, + 4.238065768732e-05, + 4.344489527284e-05, + 4.448568128282e-05, + 4.550220837700e-05,  \
+ 4.649413924199e-05, + 4.746105085360e-05, + 4.840281879297e-05, + 4.931903386023e-05, + 5.020967393648e-05,  \
+ 5.107468372444e-05, + 5.191398580791e-05, + 5.272779031657e-05, + 5.351595900720e-05, + 5.427893425804e-05,  \
+ 5.501678795554e-05, + 5.572974128881e-05, + 5.641823663609e-05, + 5.708257260267e-05, + 5.772306438303e-05 ]

* Data table for Id-Vg at Vd = 0.39V
.param vg_data_vd0.39=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.39=[ \
+ 4.020820000000e-10, + 5.842690000000e-10, + 8.489820000000e-10, + 1.233600000000e-09, + 1.792300000000e-09,  \
+ 2.603800000000e-09, + 3.782400000000e-09, + 5.493300000000e-09, + 7.976200000000e-09, + 1.157680000000e-08,  \
+ 1.679370000000e-08, + 2.434230000000e-08, + 3.524390000000e-08, + 5.094560000000e-08, + 7.347420000000e-08,  \
+ 1.056260000000e-07, + 1.511780000000e-07, + 2.150820000000e-07, + 3.035930000000e-07, + 4.242300000000e-07,  \
+ 5.854940000000e-07, + 7.963240000000e-07, + 1.065300000000e-06, + 1.400000000000e-06, + 1.806000000000e-06,  \
+ 2.286800000000e-06, + 2.843800000000e-06, + 3.476200000000e-06, + 4.181500000000e-06, + 4.956100000000e-06,  \
+ 5.795500000000e-06, + 6.694800000000e-06, + 7.648900000000e-06, + 8.652800000000e-06, + 9.701600000000e-06,  \
+ 1.079060000000e-05, + 1.191540000000e-05, + 1.307200000000e-05, + 1.425650000000e-05, + 1.546520000000e-05,  \
+ 1.669480000000e-05, + 1.794200000000e-05, + 1.920390000000e-05, + 2.047760000000e-05, + 2.176030000000e-05,  \
+ 2.304930000000e-05, + 2.434210000000e-05, + 2.563640000000e-05, + 2.692960000000e-05, + 2.821970000000e-05,  \
+ 2.950430000000e-05, + 3.078130000000e-05, + 3.204890000000e-05, + 3.330490000000e-05, + 3.454760000000e-05,  \
+ 3.577530000000e-05, + 3.698610000000e-05, + 3.817870000000e-05, + 3.935150000000e-05, + 4.050320000000e-05,  \
+ 4.163250000000e-05, + 4.273830000000e-05, + 4.381970000000e-05, + 4.487570000000e-05, + 4.590560000000e-05,  \
+ 4.690880000000e-05, + 4.788470000000e-05, + 4.883280000000e-05, + 4.975300000000e-05, + 5.064510000000e-05,  \
+ 5.150880000000e-05, + 5.234430000000e-05, + 5.315160000000e-05, + 5.393090000000e-05, + 5.468240000000e-05,  \
+ 5.540650000000e-05, + 5.610350000000e-05, + 5.677370000000e-05, + 5.741770000000e-05, + 5.803600000000e-05 ]

.param id_pred_data_vd0.39=[ \
+ 4.051814217476e-10, + 5.806258840391e-10, + 8.426942410544e-10, + 1.228111712326e-09, + 1.787723742375e-09,  \
+ 2.595146431084e-09, + 3.760922133722e-09, + 5.452283584617e-09, + 7.918256663686e-09, + 1.152068755061e-08,  \
+ 1.677343895778e-08, + 2.439711067836e-08, + 3.540049448247e-08, + 5.120273740999e-08, + 7.380447485161e-08,  \
+ 1.060009876142e-07, + 1.516109298905e-07, + 2.156669876285e-07, + 3.044961744081e-07, + 4.256183808593e-07,  \
+ 5.874116459381e-07, + 7.985644401742e-07, + 1.067383152531e-06, + 1.401107269885e-06, + 1.805325314308e-06,  \
+ 2.283658182023e-06, + 2.837641382030e-06, + 3.466871085038e-06, + 4.169316971456e-06, + 4.941638626406e-06,  \
+ 5.779609055026e-06, + 6.678459631075e-06, + 7.633116329089e-06, + 8.638497674838e-06, + 9.689571143099e-06,  \
+ 1.078152483387e-05, + 1.190975257487e-05, + 1.306994188781e-05, + 1.425800943252e-05, + 1.547013434902e-05,  \
+ 1.670278237725e-05, + 1.795246465917e-05, + 1.921607825352e-05, + 2.049055285170e-05, + 2.177304941142e-05,  \
+ 2.306080976268e-05, + 2.435130983940e-05, + 2.564198301116e-05, + 2.693057336728e-05, + 2.821484486049e-05,  \
+ 2.949263805931e-05, + 3.076204608078e-05, + 3.202113082807e-05, + 3.326823512907e-05, + 3.450163654634e-05,  \
+ 3.571987086616e-05, + 3.692163561936e-05, + 3.810546375462e-05, + 3.927035642846e-05, + 4.041528074595e-05,  \
+ 4.153907895670e-05, + 4.264106719347e-05, + 4.372043105832e-05, + 4.477674207010e-05, + 4.580918015563e-05,  \
+ 4.681744736445e-05, + 4.780106697581e-05, + 4.875980346696e-05, + 4.969344401616e-05, + 5.060189214419e-05,  \
+ 5.148490381544e-05, + 5.234257550910e-05, + 5.317486182321e-05, + 5.398196706665e-05, + 5.476401609485e-05,  \
+ 5.552111673751e-05, + 5.625358113321e-05, + 5.696164196706e-05, + 5.764562272816e-05, + 5.830600013724e-05 ]

* Data table for Id-Vg at Vd = 0.40V
.param vg_data_vd0.40=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.40=[ \
+ 4.061030000000e-10, + 5.900360000000e-10, + 8.572510000000e-10, + 1.245400000000e-09, + 1.809300000000e-09,  \
+ 2.628200000000e-09, + 3.817200000000e-09, + 5.543300000000e-09, + 8.047600000000e-09, + 1.167890000000e-08,  \
+ 1.693940000000e-08, + 2.455000000000e-08, + 3.553950000000e-08, + 5.136480000000e-08, + 7.406650000000e-08,  \
+ 1.064590000000e-07, + 1.523390000000e-07, + 2.166870000000e-07, + 3.057850000000e-07, + 4.271790000000e-07,  \
+ 5.893960000000e-07, + 8.013860000000e-07, + 1.071800000000e-06, + 1.408000000000e-06, + 1.815800000000e-06,  \
+ 2.298600000000e-06, + 2.857600000000e-06, + 3.492200000000e-06, + 4.199800000000e-06, + 4.976800000000e-06,  \
+ 5.818800000000e-06, + 6.720700000000e-06, + 7.677600000000e-06, + 8.684400000000e-06, + 9.736100000000e-06,  \
+ 1.082830000000e-05, + 1.195650000000e-05, + 1.311660000000e-05, + 1.430480000000e-05, + 1.551750000000e-05,  \
+ 1.675140000000e-05, + 1.800340000000e-05, + 1.927030000000e-05, + 2.054940000000e-05, + 2.183790000000e-05,  \
+ 2.313320000000e-05, + 2.443290000000e-05, + 2.573450000000e-05, + 2.703570000000e-05, + 2.833430000000e-05,  \
+ 2.962810000000e-05, + 3.091510000000e-05, + 3.219310000000e-05, + 3.346040000000e-05, + 3.471510000000e-05,  \
+ 3.595540000000e-05, + 3.717960000000e-05, + 3.838620000000e-05, + 3.957370000000e-05, + 4.074070000000e-05,  \
+ 4.188590000000e-05, + 4.300820000000e-05, + 4.410660000000e-05, + 4.518000000000e-05, + 4.622760000000e-05,  \
+ 4.724880000000e-05, + 4.824290000000e-05, + 4.920950000000e-05, + 5.014820000000e-05, + 5.105870000000e-05,  \
+ 5.194080000000e-05, + 5.279450000000e-05, + 5.361980000000e-05, + 5.441680000000e-05, + 5.518570000000e-05,  \
+ 5.592670000000e-05, + 5.664020000000e-05, + 5.732650000000e-05, + 5.798600000000e-05, + 5.861910000000e-05 ]

.param id_pred_data_vd0.40=[ \
+ 4.091013305896e-10, + 5.861615193226e-10, + 8.507754500897e-10, + 1.240035629735e-09, + 1.805149807410e-09,  \
+ 2.620133088271e-09, + 3.796047209903e-09, + 5.500958977223e-09, + 7.985381955677e-09, + 1.161361069535e-08,  \
+ 1.690331288273e-08, + 2.458057508647e-08, + 3.566180453163e-08, + 5.157660893929e-08, + 7.433940822921e-08,  \
+ 1.067638891072e-07, + 1.526915980321e-07, + 2.171833330067e-07, + 3.065967121074e-07, + 4.284829628887e-07,  \
+ 5.912466804148e-07, + 8.035887731239e-07, + 1.073826388165e-06, + 1.409179185430e-06, + 1.815220639401e-06,  \
+ 2.295529338880e-06, + 2.851611498045e-06, + 3.483028558549e-06, + 4.187705781078e-06, + 4.962293314748e-06,  \
+ 5.802559826407e-06, + 6.703732651658e-06, + 7.660759729333e-06, + 8.668592636241e-06, + 9.722205140861e-06,  \
+ 1.081685695681e-05, + 1.194796059281e-05, + 1.311125961365e-05, + 1.430275588064e-05, + 1.551863970235e-05,  \
+ 1.675536041148e-05, + 1.800957834348e-05, + 1.927813136717e-05, + 2.055801451206e-05, + 2.184640034102e-05,  \
+ 2.314057492185e-05, + 2.443791599944e-05, + 2.573597594164e-05, + 2.703243517317e-05, + 2.832504687831e-05,  \
+ 2.961173013318e-05, + 3.089044475928e-05, + 3.215938631911e-05, + 3.341675328556e-05, + 3.466091293376e-05,  \
+ 3.589031693991e-05, + 3.710358578246e-05, + 3.829941852018e-05, + 3.947679069825e-05, + 4.063439846504e-05,  \
+ 4.177145892754e-05, + 4.288709606044e-05, + 4.398061428219e-05, + 4.505115794018e-05, + 4.609840980265e-05,  \
+ 4.712171503343e-05, + 4.812085826416e-05, + 4.909542039968e-05, + 5.004536360502e-05, + 5.097026005387e-05,  \
+ 5.187008646317e-05, + 5.274498835206e-05, + 5.359476199374e-05, + 5.441960529424e-05, + 5.521962884814e-05,  \
+ 5.599504220299e-05, + 5.674599087797e-05, + 5.747263785452e-05, + 5.817556520924e-05, + 5.885475547984e-05 ]

* Data table for Id-Vg at Vd = 0.41V
.param vg_data_vd0.41=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.41=[ \
+ 4.101500000000e-10, + 5.958400000000e-10, + 8.655730000000e-10, + 1.257400000000e-09, + 1.826400000000e-09,  \
+ 2.652700000000e-09, + 3.852300000000e-09, + 5.593400000000e-09, + 8.119400000000e-09, + 1.178150000000e-08,  \
+ 1.708580000000e-08, + 2.475870000000e-08, + 3.583620000000e-08, + 5.178560000000e-08, + 7.466090000000e-08,  \
+ 1.072940000000e-07, + 1.535040000000e-07, + 2.182960000000e-07, + 3.079810000000e-07, + 4.301330000000e-07,  \
+ 5.933000000000e-07, + 8.064470000000e-07, + 1.078200000000e-06, + 1.416000000000e-06, + 1.825500000000e-06,  \
+ 2.310200000000e-06, + 2.871300000000e-06, + 3.508100000000e-06, + 4.218000000000e-06, + 4.997400000000e-06,  \
+ 5.841800000000e-06, + 6.746400000000e-06, + 7.705900000000e-06, + 8.715400000000e-06, + 9.770100000000e-06,  \
+ 1.086530000000e-05, + 1.199670000000e-05, + 1.316020000000e-05, + 1.435200000000e-05, + 1.556860000000e-05,  \
+ 1.680660000000e-05, + 1.806300000000e-05, + 1.933460000000e-05, + 2.061880000000e-05, + 2.191280000000e-05,  \
+ 2.321410000000e-05, + 2.452010000000e-05, + 2.582860000000e-05, + 2.713720000000e-05, + 2.844380000000e-05,  \
+ 2.974620000000e-05, + 3.104230000000e-05, + 3.233020000000e-05, + 3.360790000000e-05, + 3.487370000000e-05,  \
+ 3.612570000000e-05, + 3.736240000000e-05, + 3.858210000000e-05, + 3.978330000000e-05, + 4.096460000000e-05,  \
+ 4.212480000000e-05, + 4.326260000000e-05, + 4.437690000000e-05, + 4.546670000000e-05, + 4.653120000000e-05,  \
+ 4.756950000000e-05, + 4.858100000000e-05, + 4.956510000000e-05, + 5.052150000000e-05, + 5.144970000000e-05,  \
+ 5.234950000000e-05, + 5.322080000000e-05, + 5.406350000000e-05, + 5.487770000000e-05, + 5.566350000000e-05,  \
+ 5.642100000000e-05, + 5.715060000000e-05, + 5.785250000000e-05, + 5.852720000000e-05, + 5.917500000000e-05 ]

.param id_pred_data_vd0.41=[ \
+ 4.130719388762e-10, + 5.917750001139e-10, + 8.589771094414e-10, + 1.252135515273e-09, + 1.822843982424e-09,  \
+ 2.645527859002e-09, + 3.831764763262e-09, + 5.550462764958e-09, + 8.053632960525e-09, + 1.170786905647e-08,  \
+ 1.703458920588e-08, + 2.476523725647e-08, + 3.592396190299e-08, + 5.195045574169e-08, + 7.487281877161e-08,  \
+ 1.075224699321e-07, + 1.537640471838e-07, + 2.186847467556e-07, + 3.086741804736e-07, + 4.313118495247e-07,  \
+ 5.950298861990e-07, + 8.085486456366e-07, + 1.080186341369e-06, + 1.417159055563e-06, + 1.825014128372e-06,  \
+ 2.307302338522e-06, + 2.865495866899e-06, + 3.499116292005e-06, + 4.206065532344e-06, + 4.982969840057e-06,  \
+ 5.825570779052e-06, + 6.729110609740e-06, + 7.688558634982e-06, + 8.698845376784e-06, + 9.755037463037e-06,  \
+ 1.085236111976e-05, + 1.198633119202e-05, + 1.315268924373e-05, + 1.434748410247e-05, + 1.556697789056e-05,  \
+ 1.680764751654e-05, + 1.806619362469e-05, + 1.933945259225e-05, + 2.062448900688e-05, + 2.191844054323e-05,  \
+ 2.321865369595e-05, + 2.452247645124e-05, + 2.582751483715e-05, + 2.713143454457e-05, + 2.843195346941e-05,  \
+ 2.972692076582e-05, + 3.101442722254e-05, + 3.229255467886e-05, + 3.355954606377e-05, + 3.481370396912e-05,  \
+ 3.605350997532e-05, + 3.727762763447e-05, + 3.848472049867e-05, + 3.967357741203e-05, + 4.084311251063e-05,  \
+ 4.199246068310e-05, + 4.312066135753e-05, + 4.422713580425e-05, + 4.531106962531e-05, + 4.637196761905e-05,  \
+ 4.740939126350e-05, + 4.842289905355e-05, + 4.941215687722e-05, + 5.037711103796e-05, + 5.131739162607e-05,  \
+ 5.223295986070e-05, + 5.312380977557e-05, + 5.398998313467e-05, + 5.483146800543e-05, + 5.564843144384e-05,  \
+ 5.644095101161e-05, + 5.720922359615e-05, + 5.795363103971e-05, + 5.867430460057e-05, + 5.937148293015e-05 ]

* Data table for Id-Vg at Vd = 0.42V
.param vg_data_vd0.42=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.42=[ \
+ 4.142250000000e-10, + 6.016820000000e-10, + 8.739470000000e-10, + 1.269400000000e-09, + 1.843600000000e-09,  \
+ 2.677300000000e-09, + 3.887600000000e-09, + 5.643900000000e-09, + 8.191500000000e-09, + 1.188450000000e-08,  \
+ 1.723290000000e-08, + 2.496830000000e-08, + 3.613430000000e-08, + 5.220810000000e-08, + 7.525750000000e-08,  \
+ 1.081320000000e-07, + 1.546720000000e-07, + 2.199090000000e-07, + 3.101820000000e-07, + 4.330910000000e-07,  \
+ 5.972070000000e-07, + 8.115090000000e-07, + 1.084600000000e-06, + 1.424000000000e-06, + 1.835200000000e-06,  \
+ 2.321900000000e-06, + 2.885000000000e-06, + 3.523900000000e-06, + 4.236100000000e-06, + 5.017800000000e-06,  \
+ 5.864700000000e-06, + 6.771700000000e-06, + 7.733900000000e-06, + 8.746100000000e-06, + 9.803600000000e-06,  \
+ 1.090180000000e-05, + 1.203630000000e-05, + 1.320300000000e-05, + 1.439830000000e-05, + 1.561850000000e-05,  \
+ 1.686050000000e-05, + 1.812100000000e-05, + 1.939710000000e-05, + 2.068610000000e-05, + 2.198530000000e-05,  \
+ 2.329210000000e-05, + 2.460410000000e-05, + 2.591900000000e-05, + 2.723460000000e-05, + 2.854860000000e-05,  \
+ 2.985890000000e-05, + 3.116360000000e-05, + 3.246060000000e-05, + 3.374810000000e-05, + 3.502420000000e-05,  \
+ 3.628730000000e-05, + 3.753550000000e-05, + 3.876740000000e-05, + 3.998150000000e-05, + 4.117630000000e-05,  \
+ 4.235040000000e-05, + 4.350270000000e-05, + 4.463200000000e-05, + 4.573730000000e-05, + 4.681770000000e-05,  \
+ 4.787220000000e-05, + 4.890020000000e-05, + 4.990110000000e-05, + 5.087440000000e-05, + 5.181950000000e-05,  \
+ 5.273640000000e-05, + 5.362460000000e-05, + 5.448410000000e-05, + 5.531490000000e-05, + 5.611710000000e-05,  \
+ 5.689070000000e-05, + 5.763600000000e-05, + 5.835320000000e-05, + 5.904280000000e-05, + 5.970500000000e-05 ]

.param id_pred_data_vd0.42=[ \
+ 4.170938128212e-10, + 5.974638983552e-10, + 8.672909324048e-10, + 1.264404061452e-09, + 1.840802816844e-09,  \
+ 2.671321830405e-09, + 3.868083933156e-09, + 5.600850236931e-09, + 8.123009571648e-09, + 1.180356772323e-08,  \
+ 1.716750645642e-08, + 2.495176673278e-08, + 3.618770136882e-08, + 5.232536580024e-08, + 7.540618327084e-08,  \
+ 1.082792215357e-07, + 1.548310450517e-07, + 2.201762015375e-07, + 3.107337329311e-07, + 4.341130625107e-07,  \
+ 5.987733334223e-07, + 8.134537574733e-07, + 1.086475222110e-06, + 1.425054956599e-06, + 1.834720515035e-06,  \
+ 2.318989909327e-06, + 2.879305238821e-06, + 3.515150820022e-06, + 4.224405092828e-06, + 5.003656715417e-06,  \
+ 5.848651107954e-06, + 6.754605019523e-06, + 7.716495310888e-06, + 8.729287001188e-06, + 9.788045572350e-06,  \
+ 1.088805423933e-05, + 1.202484832902e-05, + 1.319422444794e-05, + 1.439227104129e-05, + 1.561528893944e-05,  \
+ 1.685977607849e-05, + 1.812246722693e-05, + 1.940024689247e-05, + 2.069019210467e-05, + 2.198950365710e-05,  \
+ 2.329544346139e-05, + 2.460545372742e-05, + 2.591708514956e-05, + 2.722804274526e-05, + 2.853596888599e-05,  \
+ 2.983885889989e-05, + 3.113468672382e-05, + 3.242148435675e-05, + 3.369751604623e-05, + 3.496113160509e-05,  \
+ 3.621078169090e-05, + 3.744502391783e-05, + 3.866255341563e-05, + 3.986218755017e-05, + 4.104287509108e-05,  \
+ 4.220360147883e-05, + 4.334363329690e-05, + 4.446214545169e-05, + 4.555844425340e-05, + 4.663207131671e-05,  \
+ 4.768245518790e-05, + 4.870927805314e-05, + 4.971220681909e-05, + 5.069104896393e-05, + 5.164560279809e-05,  \
+ 5.257584998617e-05, + 5.348157661501e-05, + 5.436291714432e-05, + 5.521990213310e-05, + 5.605264770566e-05,  \
+ 5.686122720363e-05, + 5.764589121100e-05, + 5.840689031174e-05, + 5.914442619542e-05, + 5.985878000502e-05 ]

* Data table for Id-Vg at Vd = 0.43V
.param vg_data_vd0.43=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.43=[ \
+ 4.183270000000e-10, + 6.075620000000e-10, + 8.823750000000e-10, + 1.281400000000e-09, + 1.860900000000e-09,  \
+ 2.702100000000e-09, + 3.923000000000e-09, + 5.694600000000e-09, + 8.264000000000e-09, + 1.198810000000e-08,  \
+ 1.738080000000e-08, + 2.517890000000e-08, + 3.643360000000e-08, + 5.263240000000e-08, + 7.585650000000e-08,  \
+ 1.089720000000e-07, + 1.558440000000e-07, + 2.215270000000e-07, + 3.123880000000e-07, + 4.360540000000e-07,  \
+ 6.011180000000e-07, + 8.165730000000e-07, + 1.091000000000e-06, + 1.432000000000e-06, + 1.845000000000e-06,  \
+ 2.333500000000e-06, + 2.898600000000e-06, + 3.539700000000e-06, + 4.254100000000e-06, + 5.038100000000e-06,  \
+ 5.887400000000e-06, + 6.796900000000e-06, + 7.761600000000e-06, + 8.776500000000e-06, + 9.836700000000e-06,  \
+ 1.093770000000e-05, + 1.207520000000e-05, + 1.324510000000e-05, + 1.444360000000e-05, + 1.566740000000e-05,  \
+ 1.691310000000e-05, + 1.817750000000e-05, + 1.945790000000e-05, + 2.075140000000e-05, + 2.205550000000e-05,  \
+ 2.336750000000e-05, + 2.468520000000e-05, + 2.600620000000e-05, + 2.732820000000e-05, + 2.864920000000e-05,  \
+ 2.996700000000e-05, + 3.127960000000e-05, + 3.258510000000e-05, + 3.388170000000e-05, + 3.516750000000e-05,  \
+ 3.644080000000e-05, + 3.769990000000e-05, + 3.894320000000e-05, + 4.016920000000e-05, + 4.137660000000e-05,  \
+ 4.256390000000e-05, + 4.372980000000e-05, + 4.487330000000e-05, + 4.599310000000e-05, + 4.708850000000e-05,  \
+ 4.815840000000e-05, + 4.920210000000e-05, + 5.021890000000e-05, + 5.120820000000e-05, + 5.216960000000e-05,  \
+ 5.310270000000e-05, + 5.400720000000e-05, + 5.488300000000e-05, + 5.572980000000e-05, + 5.654780000000e-05,  \
+ 5.733710000000e-05, + 5.809770000000e-05, + 5.882980000000e-05, + 5.953390000000e-05, + 6.021020000000e-05 ]

.param id_pred_data_vd0.43=[ \
+ 4.211650606045e-10, + 6.032243793364e-10, + 8.757098335366e-10, + 1.276840879694e-09, + 1.859015537065e-09,  \
+ 2.697520189443e-09, + 3.905006042970e-09, + 5.652090955266e-09, + 8.193588616479e-09, + 1.190079082392e-08,  \
+ 1.730227719321e-08, + 2.514030821743e-08, + 3.645356294157e-08, + 5.270225258869e-08, + 7.594098065056e-08,  \
+ 1.090363559797e-07, + 1.558962787840e-07, + 2.216622647211e-07, + 3.127811902459e-07, + 4.368943473310e-07,  \
+ 6.024859578702e-07, + 8.183133172679e-07, + 1.092710447210e-06, + 1.432883389043e-06, + 1.844349048952e-06,  \
+ 2.330601946596e-06, + 2.893046948884e-06, + 3.531142601787e-06, + 4.242716831868e-06, + 5.024359006711e-06,  \
+ 5.871774646948e-06, + 6.780190979043e-06, + 7.744580634608e-06, + 8.759889260546e-06, + 9.821254134295e-06,  \
+ 1.092396270906e-05, + 1.206358636409e-05, + 1.323593347479e-05, + 1.443716126232e-05, + 1.566360606375e-05,  \
+ 1.691178254987e-05, + 1.817849009967e-05, + 1.946066575329e-05, + 2.075534041069e-05, + 2.205973112723e-05,  \
+ 2.337117854040e-05, + 2.468707334629e-05, + 2.600506435556e-05, + 2.732271277637e-05, + 2.863778005121e-05,  \
+ 2.994820439199e-05, + 3.125188020931e-05, + 3.254690527683e-05, + 3.383154944459e-05, + 3.510414200719e-05,  \
+ 3.636299661594e-05, + 3.760676481761e-05, + 3.883414508891e-05, + 4.004391412309e-05, + 4.123502068978e-05,  \
+ 4.240651993314e-05, + 4.355747325462e-05, + 4.468725805054e-05, + 4.579504522553e-05, + 4.688037173764e-05,  \
+ 4.794288404810e-05, + 4.898209095700e-05, + 4.999769211281e-05, + 5.098939967866e-05, + 5.195720739721e-05,  \
+ 5.290088374750e-05, + 5.382052258938e-05, + 5.471600816236e-05, + 5.558735923842e-05, + 5.643473850796e-05,  \
+ 5.725838374929e-05, + 5.805838256492e-05, + 5.883481630008e-05, + 5.958826688584e-05, + 6.031862169039e-05 ]

* Data table for Id-Vg at Vd = 0.44V
.param vg_data_vd0.44=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.44=[ \
+ 4.224580000000e-10, + 6.134830000000e-10, + 8.908590000000e-10, + 1.293600000000e-09, + 1.878300000000e-09,  \
+ 2.727000000000e-09, + 3.958700000000e-09, + 5.745600000000e-09, + 8.336900000000e-09, + 1.209230000000e-08,  \
+ 1.752930000000e-08, + 2.539050000000e-08, + 3.673430000000e-08, + 5.305850000000e-08, + 7.645780000000e-08,  \
+ 1.098160000000e-07, + 1.570190000000e-07, + 2.231490000000e-07, + 3.145990000000e-07, + 4.390220000000e-07,  \
+ 6.050340000000e-07, + 8.216400000000e-07, + 1.097500000000e-06, + 1.439900000000e-06, + 1.854600000000e-06,  \
+ 2.345000000000e-06, + 2.912200000000e-06, + 3.555300000000e-06, + 4.271900000000e-06, + 5.058300000000e-06,  \
+ 5.909900000000e-06, + 6.821800000000e-06, + 7.789000000000e-06, + 8.806500000000e-06, + 9.869400000000e-06,  \
+ 1.097310000000e-05, + 1.211350000000e-05, + 1.328640000000e-05, + 1.448820000000e-05, + 1.571530000000e-05,  \
+ 1.696450000000e-05, + 1.823280000000e-05, + 1.951720000000e-05, + 2.081500000000e-05, + 2.212370000000e-05,  \
+ 2.344070000000e-05, + 2.476360000000e-05, + 2.609030000000e-05, + 2.741840000000e-05, + 2.874590000000e-05,  \
+ 3.007070000000e-05, + 3.139080000000e-05, + 3.270430000000e-05, + 3.400930000000e-05, + 3.530410000000e-05,  \
+ 3.658700000000e-05, + 3.785620000000e-05, + 3.911020000000e-05, + 4.034750000000e-05, + 4.156660000000e-05,  \
+ 4.276620000000e-05, + 4.394490000000e-05, + 4.510170000000e-05, + 4.623530000000e-05, + 4.734480000000e-05,  \
+ 4.842920000000e-05, + 4.948770000000e-05, + 5.051970000000e-05, + 5.152430000000e-05, + 5.250120000000e-05,  \
+ 5.344990000000e-05, + 5.437000000000e-05, + 5.526130000000e-05, + 5.612370000000e-05, + 5.695710000000e-05,  \
+ 5.776140000000e-05, + 5.853690000000e-05, + 5.928360000000e-05, + 6.000180000000e-05, + 6.069180000000e-05 ]

.param id_pred_data_vd0.44=[ \
+ 4.252828578188e-10, + 6.090571247341e-10, + 8.842345700089e-10, + 1.289432924878e-09, + 1.877474176126e-09,  \
+ 2.724101815232e-09, + 3.942523818523e-09, + 5.704239569582e-09, + 8.265401660879e-09, + 1.199964785314e-08,  \
+ 1.743914879171e-08, + 2.533125893933e-08, + 3.672217872008e-08, + 5.308199206411e-08, + 7.647875463590e-08,  \
+ 1.097954964280e-07, + 1.569626749642e-07, + 2.231468215541e-07, + 3.148240489281e-07, + 4.396639496917e-07,  \
+ 6.061769272492e-07, + 8.231420042648e-07, + 1.098901484511e-06, + 1.440659716536e-06, + 1.853918092820e-06,  \
+ 2.342153256905e-06, + 2.906731515395e-06, + 3.547084415914e-06, + 4.261017384124e-06, + 5.045078687544e-06,  \
+ 5.894954410905e-06, + 6.805872835685e-06, + 7.772780518280e-06, + 8.790671636234e-06, + 9.854647214524e-06,  \
+ 1.096006039006e-05, + 1.210250280565e-05, + 1.327782221779e-05, + 1.448220253224e-05, + 1.571197892190e-05,  \
+ 1.696380029898e-05, + 1.823440281441e-05, + 1.952078353497e-05, + 2.081999395159e-05, + 2.212931285612e-05,  \
+ 2.344603824895e-05, + 2.476763620507e-05, + 2.609166884213e-05, + 2.741577191046e-05, + 2.873764518881e-05,  \
+ 3.005522215972e-05, + 3.136642830214e-05, + 3.266934276326e-05, + 3.396218875423e-05, + 3.524322470184e-05,  \
+ 3.651092993096e-05, + 3.776375815505e-05, + 3.900053765392e-05, + 4.021986300359e-05, + 4.142082500039e-05,  \
+ 4.260235436959e-05, + 4.376363154734e-05, + 4.490381776122e-05, + 4.602241358953e-05, + 4.711883637356e-05,  \
+ 4.819254507311e-05, + 4.924317472614e-05, + 5.027046921896e-05, + 5.127418844495e-05, + 5.225432600128e-05,  \
+ 5.321045609890e-05, + 5.414280924015e-05, + 5.505136621650e-05, + 5.593621986918e-05, + 5.679721012712e-05,  \
+ 5.763471475802e-05, + 5.844894505572e-05, + 5.923997785430e-05, + 6.000806286465e-05, + 6.075341138057e-05 ]

* Data table for Id-Vg at Vd = 0.45V
.param vg_data_vd0.45=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.45=[ \
+ 4.266170000000e-10, + 6.194430000000e-10, + 8.993990000000e-10, + 1.305800000000e-09, + 1.895800000000e-09,  \
+ 2.752100000000e-09, + 3.994600000000e-09, + 5.796900000000e-09, + 8.410300000000e-09, + 1.219700000000e-08,  \
+ 1.767860000000e-08, + 2.560310000000e-08, + 3.703640000000e-08, + 5.348650000000e-08, + 7.706170000000e-08,  \
+ 1.106640000000e-07, + 1.581990000000e-07, + 2.247760000000e-07, + 3.168150000000e-07, + 4.419960000000e-07,  \
+ 6.089560000000e-07, + 8.267100000000e-07, + 1.103900000000e-06, + 1.447900000000e-06, + 1.864300000000e-06,  \
+ 2.356600000000e-06, + 2.925700000000e-06, + 3.571000000000e-06, + 4.289700000000e-06, + 5.078300000000e-06,  \
+ 5.932200000000e-06, + 6.846500000000e-06, + 7.816200000000e-06, + 8.836100000000e-06, + 9.901600000000e-06,  \
+ 1.100810000000e-05, + 1.215130000000e-05, + 1.332710000000e-05, + 1.453200000000e-05, + 1.576230000000e-05,  \
+ 1.701490000000e-05, + 1.828680000000e-05, + 1.957510000000e-05, + 2.087700000000e-05, + 2.219000000000e-05,  \
+ 2.351170000000e-05, + 2.483970000000e-05, + 2.617160000000e-05, + 2.750550000000e-05, + 2.883910000000e-05,  \
+ 3.017040000000e-05, + 3.149750000000e-05, + 3.281850000000e-05, + 3.413150000000e-05, + 3.543480000000e-05,  \
+ 3.672660000000e-05, + 3.800520000000e-05, + 3.926930000000e-05, + 4.051710000000e-05, + 4.174720000000e-05,  \
+ 4.295830000000e-05, + 4.414910000000e-05, + 4.531830000000e-05, + 4.646490000000e-05, + 4.758770000000e-05,  \
+ 4.868590000000e-05, + 4.975850000000e-05, + 5.080470000000e-05, + 5.182400000000e-05, + 5.281560000000e-05,  \
+ 5.377920000000e-05, + 5.471420000000e-05, + 5.562050000000e-05, + 5.649780000000e-05, + 5.734590000000e-05,  \
+ 5.816490000000e-05, + 5.895480000000e-05, + 5.971560000000e-05, + 6.044760000000e-05, + 6.115100000000e-05 ]

.param id_pred_data_vd0.45=[ \
+ 4.294450794973e-10, + 6.149545872525e-10, + 8.928578876244e-10, + 1.302171770412e-09, + 1.896167223236e-09,  \
+ 2.751045991012e-09, + 3.980623430877e-09, + 5.757222298897e-09, + 8.338450729894e-09, + 1.210018245601e-08,  \
+ 1.757807979175e-08, + 2.552478548523e-08, + 3.699397908008e-08, + 5.346539531104e-08, + 7.702042523761e-08,  \
+ 1.105594336082e-07, + 1.580335350582e-07, + 2.246345189860e-07, + 3.168670190234e-07, + 4.424284043125e-07,  \
+ 6.098580968228e-07, + 8.279512371701e-07, + 1.105062563056e-06, + 1.448394300496e-06, + 1.863442980721e-06,  \
+ 2.353650074838e-06, + 2.920372935478e-06, + 3.563003792806e-06, + 4.279308632249e-06, + 5.065807408755e-06,  \
+ 5.918198667132e-06, + 6.831634163973e-06, + 7.801115862094e-06, + 8.821606024867e-06, + 9.888232671074e-06,  \
+ 1.099637429434e-05, + 1.214160665768e-05, + 1.331987223239e-05, + 1.452736069041e-05, + 1.576043032401e-05,  \
+ 1.701577093627e-05, + 1.829019674915e-05, + 1.958064312930e-05, + 2.088427463605e-05, + 2.219833604613e-05,  \
+ 2.352017691010e-05, + 2.484725646354e-05, + 2.617711907078e-05, + 2.750741878117e-05, + 2.883585875679e-05,  \
+ 3.016035334440e-05, + 3.147881689074e-05, + 3.278927833890e-05, + 3.408995980863e-05, + 3.537915545166e-05,  \
+ 3.665524782264e-05, + 3.791678645939e-05, + 3.916242567357e-05, + 4.039093437314e-05, + 4.160116659477e-05,  \
+ 4.279224813217e-05, + 4.396322947287e-05, + 4.511343286140e-05, + 4.624210523616e-05, + 4.734877184092e-05,  \
+ 4.843294154853e-05, + 4.949423782818e-05, + 5.053240856796e-05, + 5.154740138096e-05, + 5.253872514004e-05,  \
+ 5.350648789317e-05, + 5.445062088256e-05, + 5.537131728488e-05, + 5.626844940707e-05, + 5.714206636185e-05,  \
+ 5.799257414765e-05, + 5.881993347430e-05, + 5.962445866317e-05, + 6.040622174623e-05, + 6.116562217358e-05 ]

* Data table for Id-Vg at Vd = 0.46V
.param vg_data_vd0.46=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.46=[ \
+ 4.308060000000e-10, + 6.254450000000e-10, + 9.079960000000e-10, + 1.318100000000e-09, + 1.913400000000e-09,  \
+ 2.777300000000e-09, + 4.030600000000e-09, + 5.848500000000e-09, + 8.484000000000e-09, + 1.230220000000e-08,  \
+ 1.782870000000e-08, + 2.581680000000e-08, + 3.734000000000e-08, + 5.391640000000e-08, + 7.766800000000e-08,  \
+ 1.115140000000e-07, + 1.593830000000e-07, + 2.264080000000e-07, + 3.190380000000e-07, + 4.449770000000e-07,  \
+ 6.128840000000e-07, + 8.317840000000e-07, + 1.110300000000e-06, + 1.455800000000e-06, + 1.874000000000e-06,  \
+ 2.368100000000e-06, + 2.939200000000e-06, + 3.586500000000e-06, + 4.307400000000e-06, + 5.098200000000e-06,  \
+ 5.954400000000e-06, + 6.871000000000e-06, + 7.843100000000e-06, + 8.865500000000e-06, + 9.933600000000e-06,  \
+ 1.104270000000e-05, + 1.218850000000e-05, + 1.336720000000e-05, + 1.457500000000e-05, + 1.580850000000e-05,  \
+ 1.706440000000e-05, + 1.833970000000e-05, + 1.963170000000e-05, + 2.093750000000e-05, + 2.225470000000e-05,  \
+ 2.358080000000e-05, + 2.491350000000e-05, + 2.625050000000e-05, + 2.758970000000e-05, + 2.892910000000e-05,  \
+ 3.026660000000e-05, + 3.160030000000e-05, + 3.292820000000e-05, + 3.424870000000e-05, + 3.555990000000e-05,  \
+ 3.686010000000e-05, + 3.814760000000e-05, + 3.942100000000e-05, + 4.067870000000e-05, + 4.191920000000e-05,  \
+ 4.314110000000e-05, + 4.434320000000e-05, + 4.552420000000e-05, + 4.668290000000e-05, + 4.781840000000e-05,  \
+ 4.892950000000e-05, + 5.001540000000e-05, + 5.107520000000e-05, + 5.210830000000e-05, + 5.311400000000e-05,  \
+ 5.409170000000e-05, + 5.504110000000e-05, + 5.596170000000e-05, + 5.685330000000e-05, + 5.771570000000e-05,  \
+ 5.854880000000e-05, + 5.935260000000e-05, + 6.012710000000e-05, + 6.087250000000e-05, + 6.158900000000e-05 ]

.param id_pred_data_vd0.46=[ \
+ 4.336522274606e-10, + 6.209151726111e-10, + 9.015705559889e-10, + 1.315056721296e-09, + 1.915086711435e-09,  \
+ 2.778357330868e-09, + 4.019290678059e-09, + 5.811073968687e-09, + 8.412739234132e-09, + 1.220242047850e-08,  \
+ 1.771930115524e-08, + 2.572121488242e-08, + 3.726921534053e-08, + 5.385310942074e-08, + 7.756726802199e-08,  \
+ 1.113291119736e-07, + 1.591109497667e-07, + 2.261286613248e-07, + 3.189150561411e-07, + 4.451971085473e-07,  \
+ 6.135365015325e-07, + 8.327512728101e-07, + 1.111205269808e-06, + 1.456107906961e-06, + 1.872936609288e-06,  \
+ 2.365122199990e-06, + 2.933986197604e-06, + 3.578902724257e-06, + 4.297596278775e-06, + 5.086573492008e-06,  \
+ 5.941483759671e-06, + 6.857493262942e-06, + 7.829569040041e-06, + 8.852683567966e-06, + 9.922007629939e-06,  \
+ 1.103284128476e-05, + 1.218090630573e-05, + 1.336206838459e-05, + 1.457261743781e-05, + 1.580894044309e-05,  \
+ 1.706773815386e-05, + 1.834582930314e-05, + 1.964029368537e-05, + 2.094819770718e-05, + 2.226685377536e-05,  \
+ 2.359362952120e-05, + 2.492599465768e-05, + 2.626149922435e-05, + 2.759777191386e-05, + 2.893256358220e-05,  \
+ 3.026371879969e-05, + 3.158920429996e-05, + 3.290698849014e-05, + 3.421524394071e-05, + 3.551229383447e-05,  \
+ 3.679655506858e-05, + 3.806640437688e-05, + 3.932059669751e-05, + 4.055777986650e-05, + 4.177695984254e-05,  \
+ 4.297708903323e-05, + 4.415734074428e-05, + 4.531685815891e-05, + 4.645508903195e-05, + 4.757143760798e-05,  \
+ 4.866548551945e-05, + 4.973680770490e-05, + 5.078520000097e-05, + 5.181041473406e-05, + 5.281233476126e-05,  \
+ 5.379077600082e-05, + 5.474598277942e-05, + 5.567772750510e-05, + 5.658624781063e-05, + 5.747165414505e-05,  \
+ 5.833395989612e-05, + 5.917352653341e-05, + 5.999049462844e-05, + 6.078505830374e-05, + 6.155743845738e-05 ]

* Data table for Id-Vg at Vd = 0.47V
.param vg_data_vd0.47=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.47=[ \
+ 4.350250000000e-10, + 6.314890000000e-10, + 9.166520000000e-10, + 1.330500000000e-09, + 1.931200000000e-09,  \
+ 2.802700000000e-09, + 4.067000000000e-09, + 5.900400000000e-09, + 8.558200000000e-09, + 1.240810000000e-08,  \
+ 1.797960000000e-08, + 2.603160000000e-08, + 3.764500000000e-08, + 5.434830000000e-08, + 7.827710000000e-08,  \
+ 1.123680000000e-07, + 1.605720000000e-07, + 2.280460000000e-07, + 3.212660000000e-07, + 4.479650000000e-07,  \
+ 6.168180000000e-07, + 8.368640000000e-07, + 1.116700000000e-06, + 1.463800000000e-06, + 1.883600000000e-06,  \
+ 2.379600000000e-06, + 2.952700000000e-06, + 3.602000000000e-06, + 4.325000000000e-06, + 5.118000000000e-06,  \
+ 5.976500000000e-06, + 6.895400000000e-06, + 7.869800000000e-06, + 8.894600000000e-06, + 9.965200000000e-06,  \
+ 1.107680000000e-05, + 1.222530000000e-05, + 1.340680000000e-05, + 1.461740000000e-05, + 1.585390000000e-05,  \
+ 1.711300000000e-05, + 1.839160000000e-05, + 1.968710000000e-05, + 2.099660000000e-05, + 2.231780000000e-05,  \
+ 2.364810000000e-05, + 2.498520000000e-05, + 2.632710000000e-05, + 2.767140000000e-05, + 2.901620000000e-05,  \
+ 3.035950000000e-05, + 3.169940000000e-05, + 3.303390000000e-05, + 3.436140000000e-05, + 3.568000000000e-05,  \
+ 3.698800000000e-05, + 3.828390000000e-05, + 3.956610000000e-05, + 4.083300000000e-05, + 4.208320000000e-05,  \
+ 4.331530000000e-05, + 4.452800000000e-05, + 4.572010000000e-05, + 4.689030000000e-05, + 4.803760000000e-05,  \
+ 4.916100000000e-05, + 5.025940000000e-05, + 5.133220000000e-05, + 5.237840000000e-05, + 5.339740000000e-05,  \
+ 5.438870000000e-05, + 5.535170000000e-05, + 5.628610000000e-05, + 5.719140000000e-05, + 5.806750000000e-05,  \
+ 5.891420000000e-05, + 5.973140000000e-05, + 6.051920000000e-05, + 6.127760000000e-05, + 6.200680000000e-05 ]

.param id_pred_data_vd0.47=[ \
+ 4.379006934840e-10, + 6.269336738640e-10, + 9.103720000070e-10, + 1.328069454409e-09, + 1.934210249743e-09,  \
+ 2.806005010569e-09, + 4.058489366798e-09, + 5.865755774437e-09, + 8.488243281590e-09, + 1.230632506122e-08,  \
+ 1.786282172844e-08, + 2.592064699769e-08, + 3.754823005409e-08, + 5.424562367295e-08, + 7.812010281327e-08,  \
+ 1.121063178289e-07, + 1.601971459309e-07, + 2.276332975271e-07, + 3.209745989352e-07, + 4.479747792629e-07,  \
+ 6.172219877953e-07, + 8.375538516248e-07, + 1.117348315347e-06, + 1.463808710014e-06, + 1.882412593659e-06,  \
+ 2.376574002483e-06, + 2.947588041025e-06, + 3.594791287469e-06, + 4.315897458582e-06, + 5.107362676426e-06,  \
+ 5.964828533251e-06, + 6.883425803608e-06, + 7.858128810767e-06, + 8.883916580089e-06, + 9.955892528524e-06,  \
+ 1.106947425797e-05, + 1.222033755766e-05, + 1.340442751825e-05, + 1.461797819502e-05, + 1.585749978403e-05,  \
+ 1.711965807772e-05, + 1.840139073465e-05, + 1.969968157937e-05, + 2.101176065480e-05, + 2.233486655314e-05,  \
+ 2.366643791902e-05, + 2.500391681679e-05, + 2.634485132148e-05, + 2.768695194391e-05, + 2.902785396145e-05,  \
+ 3.036551068362e-05, + 3.169774718117e-05, + 3.302267577965e-05, + 3.433828227571e-05, + 3.564291837392e-05,  \
+ 3.693500417285e-05, + 3.821291189524e-05, + 3.947535573388e-05, + 4.072101910424e-05, + 4.194874614768e-05,  \
+ 4.315759644669e-05, + 4.434669455804e-05, + 4.551513426122e-05, + 4.666253254982e-05, + 4.778805501701e-05,  \
+ 4.889137337159e-05, + 4.997210460715e-05, + 5.103002986289e-05, + 5.206495079619e-05, + 5.307665196597e-05,  \
+ 5.406520176621e-05, + 5.503042237251e-05, + 5.597256000328e-05, + 5.689164201613e-05, + 5.778771970654e-05,  \
+ 5.866102903383e-05, + 5.951177518000e-05, + 6.034021120286e-05, + 6.114646021160e-05, + 6.193098728545e-05 ]

* Data table for Id-Vg at Vd = 0.48V
.param vg_data_vd0.48=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.48=[ \
+ 4.392740000000e-10, + 6.375740000000e-10, + 9.253670000000e-10, + 1.343000000000e-09, + 1.949000000000e-09,  \
+ 2.828200000000e-09, + 4.103500000000e-09, + 5.952700000000e-09, + 8.632800000000e-09, + 1.251450000000e-08,  \
+ 1.813140000000e-08, + 2.624750000000e-08, + 3.795160000000e-08, + 5.478230000000e-08, + 7.888880000000e-08,  \
+ 1.132250000000e-07, + 1.617640000000e-07, + 2.296890000000e-07, + 3.235020000000e-07, + 4.509590000000e-07,  \
+ 6.207590000000e-07, + 8.419500000000e-07, + 1.123200000000e-06, + 1.471800000000e-06, + 1.893300000000e-06,  \
+ 2.391000000000e-06, + 2.966100000000e-06, + 3.617400000000e-06, + 4.342600000000e-06, + 5.137800000000e-06,  \
+ 5.998400000000e-06, + 6.919600000000e-06, + 7.896300000000e-06, + 8.923500000000e-06, + 9.996400000000e-06,  \
+ 1.111060000000e-05, + 1.226170000000e-05, + 1.344580000000e-05, + 1.465920000000e-05, + 1.589860000000e-05,  \
+ 1.716070000000e-05, + 1.844260000000e-05, + 1.974140000000e-05, + 2.105450000000e-05, + 2.237940000000e-05,  \
+ 2.371370000000e-05, + 2.505520000000e-05, + 2.640150000000e-05, + 2.775070000000e-05, + 2.910060000000e-05,  \
+ 3.044940000000e-05, + 3.179510000000e-05, + 3.313580000000e-05, + 3.446990000000e-05, + 3.579550000000e-05,  \
+ 3.711090000000e-05, + 3.841470000000e-05, + 3.970510000000e-05, + 4.098070000000e-05, + 4.224000000000e-05,  \
+ 4.348170000000e-05, + 4.470440000000e-05, + 4.590690000000e-05, + 4.708790000000e-05, + 4.824640000000e-05,  \
+ 4.938130000000e-05, + 5.049170000000e-05, + 5.157660000000e-05, + 5.263530000000e-05, + 5.366700000000e-05,  \
+ 5.467120000000e-05, + 5.564720000000e-05, + 5.659460000000e-05, + 5.751310000000e-05, + 5.840230000000e-05,  \
+ 5.926210000000e-05, + 6.009230000000e-05, + 6.089290000000e-05, + 6.166400000000e-05, + 6.240550000000e-05 ]

.param id_pred_data_vd0.48=[ \
+ 4.421913235575e-10, + 6.330088453410e-10, + 9.192516614576e-10, + 1.341199791227e-09, + 1.953527046794e-09,  \
+ 2.833963463900e-09, + 4.098192505353e-09, + 5.921230012973e-09, + 8.564940117139e-09, + 1.241198077651e-08,  \
+ 1.800865845780e-08, + 2.612314972339e-08, + 3.783132569879e-08, + 5.464340233630e-08, + 7.868012289691e-08,  \
+ 1.128924282057e-07, + 1.612943106011e-07, + 2.291510008945e-07, + 3.230493530282e-07, + 4.507685480348e-07,  \
+ 6.209226012288e-07, + 8.423698636761e-07, + 1.123498841480e-06, + 1.471515461162e-06, + 1.891892025014e-06,  \
+ 2.388022548985e-06, + 2.961185600725e-06, + 3.610692729126e-06, + 4.334207478678e-06, + 5.128184129717e-06,  \
+ 5.988220655126e-06, + 6.909438525327e-06, + 7.886785897426e-06, + 8.915234939195e-06, + 9.989923273679e-06,  \
+ 1.110626268201e-05, + 1.225991029060e-05, + 1.344688644167e-05, + 1.466342713684e-05, + 1.590607396793e-05,  \
+ 1.717155799270e-05, + 1.845677266829e-05, + 1.975885767024e-05, + 2.107497886755e-05, + 2.240238420200e-05,  \
+ 2.373857132625e-05, + 2.508098899852e-05, + 2.642726583872e-05, + 2.777494140901e-05, + 2.912182593718e-05,  \
+ 3.046575933695e-05, + 3.180461120792e-05, + 3.313637687825e-05, + 3.445913898759e-05, + 3.577123163268e-05,  \
+ 3.707094001584e-05, + 3.835669602267e-05, + 3.962710266933e-05, + 4.088094807230e-05, + 4.211702733301e-05,  \
+ 4.333428572863e-05, + 4.453194444068e-05, + 4.570910241455e-05, + 4.686509608291e-05, + 4.799939808436e-05,  \
+ 4.911162424833e-05, + 5.020129261538e-05, + 5.126817617565e-05, + 5.231221555732e-05, + 5.333314882591e-05,  \
+ 5.433098296635e-05, + 5.530574591830e-05, + 5.625742720440e-05, + 5.718620144762e-05, + 5.809223977849e-05,  \
+ 5.897572031245e-05, + 5.983684910461e-05, + 6.067576585338e-05, + 6.149288965389e-05, + 6.228840211406e-05 ]

* Data table for Id-Vg at Vd = 0.49V
.param vg_data_vd0.49=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.49=[ \
+ 4.435530000000e-10, + 6.437030000000e-10, + 9.341420000000e-10, + 1.355600000000e-09, + 1.967000000000e-09,  \
+ 2.853900000000e-09, + 4.140200000000e-09, + 6.005200000000e-09, + 8.707800000000e-09, + 1.262160000000e-08,  \
+ 1.828390000000e-08, + 2.646450000000e-08, + 3.825970000000e-08, + 5.521830000000e-08, + 7.950320000000e-08,  \
+ 1.140870000000e-07, + 1.629620000000e-07, + 2.313380000000e-07, + 3.257430000000e-07, + 4.539610000000e-07,  \
+ 6.247080000000e-07, + 8.470420000000e-07, + 1.129600000000e-06, + 1.479700000000e-06, + 1.902900000000e-06,  \
+ 2.402500000000e-06, + 2.979500000000e-06, + 3.632800000000e-06, + 4.360100000000e-06, + 5.157400000000e-06,  \
+ 6.020200000000e-06, + 6.943600000000e-06, + 7.922600000000e-06, + 8.952100000000e-06, + 1.002740000000e-05,  \
+ 1.114400000000e-05, + 1.229760000000e-05, + 1.348430000000e-05, + 1.470050000000e-05, + 1.594270000000e-05,  \
+ 1.720770000000e-05, + 1.849260000000e-05, + 1.979470000000e-05, + 2.111120000000e-05, + 2.243970000000e-05,  \
+ 2.377790000000e-05, + 2.512340000000e-05, + 2.647400000000e-05, + 2.782780000000e-05, + 2.918260000000e-05,  \
+ 3.053650000000e-05, + 3.188770000000e-05, + 3.323430000000e-05, + 3.457460000000e-05, + 3.590670000000e-05,  \
+ 3.722920000000e-05, + 3.854030000000e-05, + 3.983850000000e-05, + 4.112220000000e-05, + 4.239020000000e-05,  \
+ 4.364090000000e-05, + 4.487300000000e-05, + 4.608520000000e-05, + 4.727650000000e-05, + 4.844550000000e-05,  \
+ 4.959140000000e-05, + 5.071300000000e-05, + 5.180940000000e-05, + 5.287990000000e-05, + 5.392370000000e-05,  \
+ 5.494010000000e-05, + 5.592850000000e-05, + 5.688850000000e-05, + 5.781950000000e-05, + 5.872130000000e-05,  \
+ 5.959370000000e-05, + 6.043640000000e-05, + 6.124940000000e-05, + 6.203260000000e-05, + 6.278610000000e-05 ]

.param id_pred_data_vd0.49=[ \
+ 4.465209146876e-10, + 6.391384987925e-10, + 9.282044133307e-10, + 1.354440255508e-09, + 1.973008076916e-09,  \
+ 2.862202781451e-09, + 4.138382188046e-09, + 5.977461272622e-09, + 8.642782525214e-09, + 1.251931694313e-08,  \
+ 1.815680853667e-08, + 2.632886200615e-08, + 3.811876347015e-08, + 5.504681780621e-08, + 7.924738667953e-08,  \
+ 1.136884698383e-07, + 1.624042312187e-07, + 2.306847528644e-07, + 3.251414761962e-07, + 4.535831226349e-07,  \
+ 6.246470763926e-07, + 8.472068896026e-07, + 1.129666786710e-06, + 1.479238426327e-06, + 1.901382443066e-06,  \
+ 2.399484346824e-06, + 2.974794192596e-06, + 3.626601387623e-06, + 4.352544419817e-06, + 5.149050048203e-06,  \
+ 6.011662862875e-06, + 6.935527926544e-06, + 7.915539845271e-06, + 8.946671659942e-06, + 1.002405952022e-05,  \
+ 1.114312924983e-05, + 1.229958565091e-05, + 1.348939913441e-05, + 1.470891713325e-05, + 1.595461275429e-05,  \
+ 1.722333345242e-05, + 1.851199798693e-05, + 1.981769713893e-05, + 2.113771777658e-05, + 2.246931111586e-05,  \
+ 2.381001180765e-05, + 2.515723506804e-05, + 2.650859220012e-05, + 2.786174263747e-05, + 2.921445277025e-05,  \
+ 3.056443907553e-05, + 3.190972820448e-05, + 3.324820776470e-05, + 3.457797392912e-05, + 3.589726191422e-05,  \
+ 3.720442102349e-05, + 3.849781838653e-05, + 3.977612417657e-05, + 4.103797291464e-05, + 4.228206686093e-05,  \
+ 4.350761810201e-05, + 4.471356776776e-05, + 4.589902455336e-05, + 4.706346080638e-05, + 4.820628826565e-05,  \
+ 4.932697571348e-05, + 5.042517019319e-05, + 5.150069344381e-05, + 5.255327807390e-05, + 5.358295260521e-05,  \
+ 5.458951738547e-05, + 5.557311145822e-05, + 5.653370273649e-05, + 5.747164417699e-05, + 5.838682525791e-05,  \
+ 5.927959180553e-05, + 6.015026825480e-05, + 6.099892591010e-05, + 6.182594268466e-05, + 6.263167510042e-05 ]

* Data table for Id-Vg at Vd = 0.50V
.param vg_data_vd0.50=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.50=[ \
+ 4.478640000000e-10, + 6.498760000000e-10, + 9.429780000000e-10, + 1.368200000000e-09, + 1.985100000000e-09,  \
+ 2.879800000000e-09, + 4.177200000000e-09, + 6.058000000000e-09, + 8.783200000000e-09, + 1.272920000000e-08,  \
+ 1.843730000000e-08, + 2.668270000000e-08, + 3.856930000000e-08, + 5.565640000000e-08, + 8.012050000000e-08,  \
+ 1.149510000000e-07, + 1.641640000000e-07, + 2.329930000000e-07, + 3.279920000000e-07, + 4.569710000000e-07,  \
+ 6.286650000000e-07, + 8.521420000000e-07, + 1.136000000000e-06, + 1.487700000000e-06, + 1.912500000000e-06,  \
+ 2.413900000000e-06, + 2.992800000000e-06, + 3.648200000000e-06, + 4.377500000000e-06, + 5.176900000000e-06,  \
+ 6.041900000000e-06, + 6.967500000000e-06, + 7.948700000000e-06, + 8.980500000000e-06, + 1.005820000000e-05,  \
+ 1.117720000000e-05, + 1.233320000000e-05, + 1.352240000000e-05, + 1.474120000000e-05, + 1.598610000000e-05,  \
+ 1.725400000000e-05, + 1.854190000000e-05, + 1.984700000000e-05, + 2.116680000000e-05, + 2.249880000000e-05,  \
+ 2.384060000000e-05, + 2.519000000000e-05, + 2.654470000000e-05, + 2.790280000000e-05, + 2.926230000000e-05,  \
+ 3.062110000000e-05, + 3.197750000000e-05, + 3.332970000000e-05, + 3.467580000000e-05, + 3.601410000000e-05,  \
+ 3.734320000000e-05, + 3.866120000000e-05, + 3.996670000000e-05, + 4.125820000000e-05, + 4.253420000000e-05,  \
+ 4.379330000000e-05, + 4.503430000000e-05, + 4.625580000000e-05, + 4.745670000000e-05, + 4.863570000000e-05,  \
+ 4.979180000000e-05, + 5.092410000000e-05, + 5.203150000000e-05, + 5.311320000000e-05, + 5.416840000000e-05,  \
+ 5.519640000000e-05, + 5.619670000000e-05, + 5.716850000000e-05, + 5.811160000000e-05, + 5.902550000000e-05,  \
+ 5.990990000000e-05, + 6.076460000000e-05, + 6.158950000000e-05, + 6.238450000000e-05, + 6.314960000000e-05 ]

.param id_pred_data_vd0.50=[ \
+ 4.508873829856e-10, + 6.453146905727e-10, + 9.372239651029e-10, + 1.367773783123e-09, + 1.992651599281e-09,  \
+ 2.890710115722e-09, + 4.179002033311e-09, + 6.034417410206e-09, + 8.721740663020e-09, + 1.262824600445e-08,  \
+ 1.830724372098e-08, + 2.653769293204e-08, + 3.841040907560e-08, + 5.545602732582e-08, + 7.982271910123e-08,  \
+ 1.144951653487e-07, + 1.635288384705e-07, + 2.322365588725e-07, + 3.272575099800e-07, + 4.564240612126e-07,  \
+ 6.283981974775e-07, + 8.520742653673e-07, + 1.135864522439e-06, + 1.486989503974e-06, + 1.910898845381e-06,  \
+ 2.410967454125e-06, + 2.988426103911e-06, + 3.642535830295e-06, + 4.370917849883e-06, + 5.169938049221e-06,  \
+ 6.035169008101e-06, + 6.961670806049e-06, + 7.944368917379e-06, + 8.978194273368e-06, + 1.005830381473e-05,  \
+ 1.118010914070e-05, + 1.233930925082e-05, + 1.353197149001e-05, + 1.475436692999e-05, + 1.600310315553e-05,  \
+ 1.727497146931e-05, + 1.856693415903e-05, + 1.987622272281e-05, + 2.119999953720e-05, + 2.253564525745e-05,  \
+ 2.388069151493e-05, + 2.523251532693e-05, + 2.658885387063e-05, + 2.794732790790e-05, + 2.930564733106e-05,  \
+ 3.066157296416e-05, + 3.201308936696e-05, + 3.335806832183e-05, + 3.469467992545e-05, + 3.602109791245e-05,  \
+ 3.733551056939e-05, + 3.863644815283e-05, + 3.992244091933e-05, + 4.119207005715e-05, + 4.244423689670e-05,  \
+ 4.367774090497e-05, + 4.489178536460e-05, + 4.608543895301e-05, + 4.725807593786e-05, + 4.840908877668e-05,  \
+ 4.953808092978e-05, + 5.064440847491e-05, + 5.172830788069e-05, + 5.278916796669e-05, + 5.382710878621e-05,  \
+ 5.484186840476e-05, + 5.583383972407e-05, + 5.680284084519e-05, + 5.774921373813e-05, + 5.867306390428e-05,  \
+ 5.957452958683e-05, + 6.045391273801e-05, + 6.131154077593e-05, + 6.214765744517e-05, + 6.296249921434e-05 ]

* Data table for Id-Vg at Vd = 0.51V
.param vg_data_vd0.51=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.51=[ \
+ 4.522070000000e-10, + 6.560930000000e-10, + 9.518760000000e-10, + 1.380900000000e-09, + 2.003300000000e-09,  \
+ 2.905800000000e-09, + 4.214500000000e-09, + 6.111200000000e-09, + 8.859200000000e-09, + 1.283750000000e-08,  \
+ 1.859150000000e-08, + 2.690200000000e-08, + 3.888060000000e-08, + 5.609670000000e-08, + 8.074070000000e-08,  \
+ 1.158200000000e-07, + 1.653710000000e-07, + 2.346530000000e-07, + 3.302480000000e-07, + 4.599890000000e-07,  \
+ 6.326300000000e-07, + 8.572500000000e-07, + 1.142500000000e-06, + 1.495600000000e-06, + 1.922200000000e-06,  \
+ 2.425300000000e-06, + 3.006100000000e-06, + 3.663500000000e-06, + 4.394900000000e-06, + 5.196400000000e-06,  \
+ 6.063500000000e-06, + 6.991300000000e-06, + 7.974700000000e-06, + 9.008700000000e-06, + 1.008870000000e-05,  \
+ 1.121000000000e-05, + 1.236840000000e-05, + 1.356010000000e-05, + 1.478140000000e-05, + 1.602900000000e-05,  \
+ 1.729960000000e-05, + 1.859040000000e-05, + 1.989850000000e-05, + 2.122150000000e-05, + 2.255680000000e-05,  \
+ 2.390210000000e-05, + 2.525510000000e-05, + 2.661380000000e-05, + 2.797600000000e-05, + 2.933990000000e-05,  \
+ 3.070340000000e-05, + 3.206470000000e-05, + 3.342210000000e-05, + 3.477370000000e-05, + 3.611800000000e-05,  \
+ 3.745320000000e-05, + 3.877780000000e-05, + 4.009020000000e-05, + 4.138890000000e-05, + 4.267260000000e-05,  \
+ 4.393970000000e-05, + 4.518900000000e-05, + 4.641930000000e-05, + 4.762920000000e-05, + 4.881760000000e-05,  \
+ 4.998350000000e-05, + 5.112580000000e-05, + 5.224350000000e-05, + 5.333590000000e-05, + 5.440190000000e-05,  \
+ 5.544100000000e-05, + 5.645250000000e-05, + 5.743570000000e-05, + 5.839030000000e-05, + 5.931570000000e-05,  \
+ 6.021170000000e-05, + 6.107790000000e-05, + 6.191420000000e-05, + 6.272060000000e-05, + 6.349690000000e-05 ]

.param id_pred_data_vd0.51=[ \
+ 4.552932914015e-10, + 6.515384731731e-10, + 9.463009675859e-10, + 1.381197116679e-09, + 2.012430089238e-09,  \
+ 2.919458075290e-09, + 4.220022731261e-09, + 6.092035889083e-09, + 8.801760920107e-09, + 1.273876103269e-08,  \
+ 1.845999214822e-08, + 2.674962043869e-08, + 3.870637144132e-08, + 5.587149708219e-08, + 8.040632309303e-08,  \
+ 1.153133550247e-07, + 1.646686831691e-07, + 2.338087116982e-07, + 3.293975208862e-07, + 4.592957157001e-07,  \
+ 6.321835974177e-07, + 8.569782153245e-07, + 1.142102075846e-06, + 1.494774710409e-06, + 1.920447425618e-06,  \
+ 2.422485513307e-06, + 3.002090325026e-06, + 3.658503478619e-06, + 4.389316472952e-06, + 5.190883275645e-06,  \
+ 6.058712733648e-06, + 6.987875131017e-06, + 7.973245938047e-06, + 9.009788755066e-06, + 1.009260262435e-05,  \
+ 1.121712055465e-05, + 1.237908354597e-05, + 1.357452945740e-05, + 1.479978094721e-05, + 1.605147237569e-05,  \
+ 1.732639117108e-05, + 1.862166707724e-05, + 1.993432222662e-05, + 2.126172385033e-05, + 2.260127999762e-05,  \
+ 2.395049519691e-05, + 2.530687583203e-05, + 2.666797281563e-05, + 2.803153187415e-05, + 2.939528945717e-05,  \
+ 3.075703396462e-05, + 3.211459646991e-05, + 3.346601028170e-05, + 3.480926789052e-05, + 3.614255103457e-05,  \
+ 3.746421585674e-05, + 3.877252573147e-05, + 4.006602604932e-05, + 4.134337723372e-05, + 4.260339555913e-05,  \
+ 4.384482308524e-05, + 4.506682118517e-05, + 4.626857349649e-05, + 4.744926365674e-05, + 4.860827197263e-05,  \
+ 4.974523108103e-05, + 5.085986638733e-05, + 5.195154706598e-05, + 5.302047720761e-05, + 5.406626347394e-05,  \
+ 5.508905429451e-05, + 5.608892017335e-05, + 5.706593903597e-05, + 5.802028899780e-05, + 5.895207767026e-05,  \
+ 5.986159449094e-05, + 6.074909921153e-05, + 6.161496661662e-05, + 6.245951211895e-05, + 6.328296949505e-05 ]

* Data table for Id-Vg at Vd = 0.52V
.param vg_data_vd0.52=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.52=[ \
+ 4.565820000000e-10, + 6.623550000000e-10, + 9.608370000000e-10, + 1.393800000000e-09, + 2.021600000000e-09,  \
+ 2.932100000000e-09, + 4.251900000000e-09, + 6.164700000000e-09, + 8.935500000000e-09, + 1.294640000000e-08,  \
+ 1.874670000000e-08, + 2.712260000000e-08, + 3.919350000000e-08, + 5.653920000000e-08, + 8.136380000000e-08,  \
+ 1.166920000000e-07, + 1.665830000000e-07, + 2.363200000000e-07, + 3.325120000000e-07, + 4.630160000000e-07,  \
+ 6.366050000000e-07, + 8.623660000000e-07, + 1.148900000000e-06, + 1.503600000000e-06, + 1.931800000000e-06,  \
+ 2.436800000000e-06, + 3.019400000000e-06, + 3.678800000000e-06, + 4.412200000000e-06, + 5.215700000000e-06,  \
+ 6.085000000000e-06, + 7.014900000000e-06, + 8.000500000000e-06, + 9.036700000000e-06, + 1.011890000000e-05,  \
+ 1.124250000000e-05, + 1.240330000000e-05, + 1.359740000000e-05, + 1.482120000000e-05, + 1.607130000000e-05,  \
+ 1.734460000000e-05, + 1.863810000000e-05, + 1.994920000000e-05, + 2.127520000000e-05, + 2.261370000000e-05,  \
+ 2.396230000000e-05, + 2.531890000000e-05, + 2.668130000000e-05, + 2.804750000000e-05, + 2.941550000000e-05,  \
+ 3.078350000000e-05, + 3.214950000000e-05, + 3.351180000000e-05, + 3.486870000000e-05, + 3.621850000000e-05,  \
+ 3.755960000000e-05, + 3.889040000000e-05, + 4.020930000000e-05, + 4.151490000000e-05, + 4.280570000000e-05,  \
+ 4.408040000000e-05, + 4.533760000000e-05, + 4.657610000000e-05, + 4.779460000000e-05, + 4.899190000000e-05,  \
+ 5.016700000000e-05, + 5.131880000000e-05, + 5.244640000000e-05, + 5.354870000000e-05, + 5.462510000000e-05,  \
+ 5.567470000000e-05, + 5.669690000000e-05, + 5.769090000000e-05, + 5.865640000000e-05, + 5.959290000000e-05,  \
+ 6.049990000000e-05, + 6.137720000000e-05, + 6.222450000000e-05, + 6.304180000000e-05, + 6.382890000000e-05 ]

.param id_pred_data_vd0.52=[ \
+ 4.597346925372e-10, + 6.578051348072e-10, + 9.554319557736e-10, + 1.394689395084e-09, + 2.032321031464e-09,  \
+ 2.948404400627e-09, + 4.261425061713e-09, + 6.150278686334e-09, + 8.882741511229e-09, + 1.285074226587e-08,  \
+ 1.861480811272e-08, + 2.696469991292e-08, + 3.900679985236e-08, + 5.629280764197e-08, + 8.099850617782e-08,  \
+ 1.161434630603e-07, + 1.658246708303e-07, + 2.354026810281e-07, + 3.315666367598e-07, + 4.621994116860e-07,  \
+ 6.360086672430e-07, + 8.619258233011e-07, + 1.148382552856e-06, + 1.502607583461e-06, + 1.930043299581e-06,  \
+ 2.434039633954e-06, + 3.015793354280e-06, + 3.674508625409e-06, + 4.407762353367e-06, + 5.211862553551e-06,  \
+ 6.082311592763e-06, + 7.014123293629e-06, + 8.002188042155e-06, + 9.041415614774e-06, + 1.012695793179e-05,  \
+ 1.125417737057e-05, + 1.241886573553e-05, + 1.361703616567e-05, + 1.484511893068e-05, + 1.609966158867e-05,  \
+ 1.737759856042e-05, + 1.867595317890e-05, + 1.999195781536e-05, + 2.132285240805e-05, + 2.266619470902e-05,  \
+ 2.401942139841e-05, + 2.538009212003e-05, + 2.674581759493e-05, + 2.811432204908e-05, + 2.948334484245e-05,  \
+ 3.085066884523e-05, + 3.221414313884e-05, + 3.357179841259e-05, + 3.492159914458e-05, + 3.626171033829e-05,  \
+ 3.759034996619e-05, + 3.890591760864e-05, + 4.020685824798e-05, + 4.149182874244e-05, + 4.275958810467e-05,  \
+ 4.400884616189e-05, + 4.523882351350e-05, + 4.644843807910e-05, + 4.763703153003e-05, + 4.880407417659e-05,  \
+ 4.994894552510e-05, + 5.107141099870e-05, + 5.217096739216e-05, + 5.324766010744e-05, + 5.430119024822e-05,  \
+ 5.533174698940e-05, + 5.633913737256e-05, + 5.732373974752e-05, + 5.828556924826e-05, + 5.922494747210e-05,  \
+ 6.014205981046e-05, + 6.103727326263e-05, + 6.191073160153e-05, + 6.276309693931e-05, + 6.359438062645e-05 ]

* Data table for Id-Vg at Vd = 0.53V
.param vg_data_vd0.53=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.53=[ \
+ 4.609890000000e-10, + 6.686620000000e-10, + 9.698610000000e-10, + 1.406700000000e-09, + 2.040100000000e-09,  \
+ 2.958400000000e-09, + 4.289600000000e-09, + 6.218600000000e-09, + 9.012400000000e-09, + 1.305600000000e-08,  \
+ 1.890270000000e-08, + 2.734440000000e-08, + 3.950800000000e-08, + 5.698390000000e-08, + 8.198990000000e-08,  \
+ 1.175680000000e-07, + 1.678000000000e-07, + 2.379930000000e-07, + 3.347830000000e-07, + 4.660510000000e-07,  \
+ 6.405880000000e-07, + 8.674910000000e-07, + 1.155400000000e-06, + 1.511500000000e-06, + 1.941400000000e-06,  \
+ 2.448200000000e-06, + 3.032700000000e-06, + 3.694000000000e-06, + 4.429400000000e-06, + 5.235000000000e-06,  \
+ 6.106400000000e-06, + 7.038400000000e-06, + 8.026100000000e-06, + 9.064600000000e-06, + 1.014890000000e-05,  \
+ 1.127480000000e-05, + 1.243790000000e-05, + 1.363430000000e-05, + 1.486050000000e-05, + 1.611310000000e-05,  \
+ 1.738900000000e-05, + 1.868520000000e-05, + 1.999910000000e-05, + 2.132800000000e-05, + 2.266960000000e-05,  \
+ 2.402140000000e-05, + 2.538140000000e-05, + 2.674740000000e-05, + 2.811740000000e-05, + 2.948940000000e-05,  \
+ 3.086160000000e-05, + 3.223200000000e-05, + 3.359910000000e-05, + 3.496100000000e-05, + 3.631600000000e-05,  \
+ 3.766270000000e-05, + 3.899930000000e-05, + 4.032440000000e-05, + 4.163640000000e-05, + 4.293410000000e-05,  \
+ 4.421590000000e-05, + 4.548060000000e-05, + 4.672680000000e-05, + 4.795340000000e-05, + 4.915920000000e-05,  \
+ 5.034300000000e-05, + 5.150380000000e-05, + 5.264060000000e-05, + 5.375250000000e-05, + 5.483860000000e-05,  \
+ 5.589820000000e-05, + 5.693050000000e-05, + 5.793490000000e-05, + 5.891090000000e-05, + 5.985790000000e-05,  \
+ 6.077550000000e-05, + 6.166330000000e-05, + 6.252130000000e-05, + 6.334900000000e-05, + 6.414650000000e-05 ]

.param id_pred_data_vd0.53=[ \
+ 4.642115053466e-10, + 6.641132033192e-10, + 9.646088472426e-10, + 1.408243868184e-09, + 2.052315135614e-09,  \
+ 2.977524382608e-09, + 4.303135741068e-09, + 6.209067962004e-09, + 8.964639821585e-09, + 1.296412964535e-08,  \
+ 1.877178529952e-08, + 2.718275560198e-08, + 3.931143872649e-08, + 5.672044181892e-08, + 8.159950155573e-08,  \
+ 1.169860270522e-07, + 1.669977029906e-07, + 2.370188590817e-07, + 3.337634581158e-07, + 4.651397352973e-07,  \
+ 6.398758625892e-07, + 8.669186286170e-07, + 1.154714261702e-06, + 1.510488846179e-06, + 1.939685489560e-06,  \
+ 2.445644554427e-06, + 3.029533522749e-06, + 3.690556559377e-06, + 4.426235536812e-06, + 5.232877365415e-06,  \
+ 6.105933589424e-06, + 7.040404088912e-06, + 8.031151846808e-06, + 9.073076962522e-06, + 1.016130609059e-05,  \
+ 1.129122811108e-05, + 1.245861078132e-05, + 1.365948215607e-05, + 1.489030026278e-05, + 1.614766002604e-05,  \
+ 1.742847547575e-05, + 1.872986405942e-05, + 2.004903577472e-05, + 2.138336258213e-05, + 2.273028007039e-05,  \
+ 2.408737807855e-05, + 2.545214232669e-05, + 2.682233232917e-05, + 2.819558420015e-05, + 2.956969216029e-05,  \
+ 3.094240801147e-05, + 3.231163394958e-05, + 3.367532037373e-05, + 3.503152373014e-05, + 3.637824454927e-05,  \
+ 3.771378222154e-05, + 3.903646313120e-05, + 4.034481033159e-05, + 4.163728131971e-05, + 4.291263823688e-05,  \
+ 4.416969335580e-05, + 4.540745947452e-05, + 4.662500723498e-05, + 4.782158466696e-05, + 4.899650921288e-05,  \
+ 5.014924485295e-05, + 5.127948694280e-05, + 5.238672260020e-05, + 5.347102895030e-05, + 5.453225559904e-05,  \
+ 5.557016731473e-05, + 5.658507645421e-05, + 5.757694445492e-05, + 5.854609524249e-05, + 5.949273705482e-05,  \
+ 6.041704727977e-05, + 6.131933827419e-05, + 6.220009207027e-05, + 6.305957089353e-05, + 6.389825677616e-05 ]

* Data table for Id-Vg at Vd = 0.54V
.param vg_data_vd0.54=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.54=[ \
+ 4.654290000000e-10, + 6.750150000000e-10, + 9.789500000000e-10, + 1.419700000000e-09, + 2.058700000000e-09,  \
+ 2.985000000000e-09, + 4.327600000000e-09, + 6.272800000000e-09, + 9.089700000000e-09, + 1.316620000000e-08,  \
+ 1.905960000000e-08, + 2.756740000000e-08, + 3.982430000000e-08, + 5.743090000000e-08, + 8.261900000000e-08,  \
+ 1.184490000000e-07, + 1.690220000000e-07, + 2.396730000000e-07, + 3.370620000000e-07, + 4.690950000000e-07,  \
+ 6.445810000000e-07, + 8.726250000000e-07, + 1.161800000000e-06, + 1.519500000000e-06, + 1.951000000000e-06,  \
+ 2.459600000000e-06, + 3.046000000000e-06, + 3.709200000000e-06, + 4.446600000000e-06, + 5.254300000000e-06,  \
+ 6.127700000000e-06, + 7.061800000000e-06, + 8.051600000000e-06, + 9.092200000000e-06, + 1.017880000000e-05,  \
+ 1.130680000000e-05, + 1.247210000000e-05, + 1.367090000000e-05, + 1.489940000000e-05, + 1.615450000000e-05,  \
+ 1.743280000000e-05, + 1.873170000000e-05, + 2.004830000000e-05, + 2.138000000000e-05, + 2.272450000000e-05,  \
+ 2.407950000000e-05, + 2.544270000000e-05, + 2.681220000000e-05, + 2.818580000000e-05, + 2.956160000000e-05,  \
+ 3.093780000000e-05, + 3.231250000000e-05, + 3.368400000000e-05, + 3.505060000000e-05, + 3.641070000000e-05,  \
+ 3.776260000000e-05, + 3.910480000000e-05, + 4.043570000000e-05, + 4.175390000000e-05, + 4.305800000000e-05,  \
+ 4.434660000000e-05, + 4.561830000000e-05, + 4.687190000000e-05, + 4.810610000000e-05, + 4.931980000000e-05,  \
+ 5.051190000000e-05, + 5.168120000000e-05, + 5.282680000000e-05, + 5.394780000000e-05, + 5.504320000000e-05,  \
+ 5.611230000000e-05, + 5.715420000000e-05, + 5.816850000000e-05, + 5.915440000000e-05, + 6.011140000000e-05,  \
+ 6.103910000000e-05, + 6.193710000000e-05, + 6.280520000000e-05, + 6.364300000000e-05, + 6.445060000000e-05 ]

.param id_pred_data_vd0.54=[ \
+ 4.687250687585e-10, + 6.704591681839e-10, + 9.738298767381e-10, + 1.421846760330e-09, + 2.072384583940e-09,  \
+ 3.006796172045e-09, + 4.345124580141e-09, + 6.268362628958e-09, + 9.047367655057e-09, + 1.307885096224e-08,  \
+ 1.893071235770e-08, + 2.740379507316e-08, + 3.962029680338e-08, + 5.715408050833e-08, + 8.220915788115e-08,  \
+ 1.178408462010e-07, + 1.681879621174e-07, + 2.386583372527e-07, + 3.359913716849e-07, + 4.681169116338e-07,  \
+ 6.437872571041e-07, + 8.719633297005e-07, + 1.161099207820e-06, + 1.518426861367e-06, + 1.949384418367e-06,  \
+ 2.457296932334e-06, + 3.043329234060e-06, + 3.706644565682e-06, + 4.444746773515e-06, + 5.253919989627e-06,  \
+ 6.129586909083e-06, + 7.066713478707e-06, + 8.060148757068e-06, + 9.104750643019e-06, + 1.019564126182e-05,  \
+ 1.132823545049e-05, + 1.249826433195e-05, + 1.370182049868e-05, + 1.493530005973e-05, + 1.619537906663e-05,  \
+ 1.747902824718e-05, + 1.878331459011e-05, + 2.010554082517e-05, + 2.144307647541e-05, + 2.279345018906e-05,  \
+ 2.415420633042e-05, + 2.552297373768e-05, + 2.689738910703e-05, + 2.827518539561e-05, + 2.965416235384e-05,  \
+ 3.103207061940e-05, + 3.240690246457e-05, + 3.377644781722e-05, + 3.513876770739e-05, + 3.649201156804e-05,  \
+ 3.783435633522e-05, + 3.916406931239e-05, + 4.047962604091e-05, + 4.177956492640e-05, + 4.306256581913e-05,  \
+ 4.432735178852e-05, + 4.557283842587e-05, + 4.679825957282e-05, + 4.800266833627e-05, + 4.918546750559e-05,  \
+ 5.034610701841e-05, + 5.148402502527e-05, + 5.259908793960e-05, + 5.369091071771e-05, + 5.475958372699e-05,  \
+ 5.580496159382e-05, + 5.682708753739e-05, + 5.782622873085e-05, + 5.880238124519e-05, + 5.975590262096e-05,  \
+ 6.068719361792e-05, + 6.159633674542e-05, + 6.248381134355e-05, + 6.335011246847e-05, + 6.419553872547e-05 ]

* Data table for Id-Vg at Vd = 0.55V
.param vg_data_vd0.55=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.55=[ \
+ 4.699020000000e-10, + 6.814150000000e-10, + 9.881040000000e-10, + 1.432800000000e-09, + 2.077400000000e-09,  \
+ 3.011800000000e-09, + 4.365800000000e-09, + 6.327300000000e-09, + 9.167500000000e-09, + 1.327700000000e-08,  \
+ 1.921740000000e-08, + 2.779160000000e-08, + 4.014220000000e-08, + 5.788020000000e-08, + 8.325120000000e-08,  \
+ 1.193330000000e-07, + 1.702500000000e-07, + 2.413590000000e-07, + 3.393490000000e-07, + 4.721480000000e-07,  \
+ 6.485840000000e-07, + 8.777690000000e-07, + 1.168300000000e-06, + 1.527500000000e-06, + 1.960600000000e-06,  \
+ 2.470900000000e-06, + 3.059200000000e-06, + 3.724400000000e-06, + 4.463800000000e-06, + 5.273500000000e-06,  \
+ 6.148900000000e-06, + 7.085100000000e-06, + 8.077000000000e-06, + 9.119700000000e-06, + 1.020840000000e-05,  \
+ 1.133860000000e-05, + 1.250610000000e-05, + 1.370710000000e-05, + 1.493800000000e-05, + 1.619540000000e-05,  \
+ 1.747620000000e-05, + 1.877760000000e-05, + 2.009680000000e-05, + 2.143130000000e-05, + 2.277860000000e-05,  \
+ 2.413660000000e-05, + 2.550300000000e-05, + 2.687570000000e-05, + 2.825280000000e-05, + 2.963220000000e-05,  \
+ 3.101230000000e-05, + 3.239100000000e-05, + 3.376680000000e-05, + 3.513800000000e-05, + 3.650280000000e-05,  \
+ 3.785970000000e-05, + 3.920710000000e-05, + 4.054360000000e-05, + 4.186760000000e-05, + 4.317780000000e-05,  \
+ 4.447280000000e-05, + 4.575120000000e-05, + 4.701170000000e-05, + 4.825320000000e-05, + 4.947450000000e-05,  \
+ 5.067430000000e-05, + 5.185170000000e-05, + 5.300570000000e-05, + 5.413520000000e-05, + 5.523940000000e-05,  \
+ 5.631750000000e-05, + 5.736870000000e-05, + 5.839220000000e-05, + 5.938760000000e-05, + 6.035420000000e-05,  \
+ 6.129160000000e-05, + 6.219930000000e-05, + 6.307710000000e-05, + 6.392470000000e-05, + 6.474180000000e-05 ]

.param id_pred_data_vd0.55=[ \
+ 4.732745445546e-10, + 6.768440197202e-10, + 9.830831926294e-10, + 1.435488516943e-09, + 2.092515205554e-09,  \
+ 3.036177087523e-09, + 4.387348750967e-09, + 6.328081481044e-09, + 9.130843903193e-09, + 1.319474192130e-08,  \
+ 1.909142728351e-08, + 2.762743189777e-08, + 3.993319026563e-08, + 5.759358181479e-08, + 8.282734356158e-08,  \
+ 1.187080705733e-07, + 1.693959731597e-07, + 2.403220719316e-07, + 3.382494242032e-07, + 4.711348594810e-07,  \
+ 6.477449574049e-07, + 8.770594547514e-07, + 1.167539858216e-06, + 1.526423068299e-06, + 1.959140058716e-06,  \
+ 2.469008177286e-06, + 3.057165554310e-06, + 3.722772316905e-06, + 4.463298091650e-06, + 5.274988461679e-06,  \
+ 6.153245385576e-06, + 7.093028625604e-06, + 8.089121865851e-06, + 9.136398330156e-06, + 1.022994883897e-05,  \
+ 1.136516184488e-05, + 1.253780847037e-05, + 1.374398098051e-05, + 1.498008377894e-05, + 1.624281039767e-05,  \
+ 1.752914849931e-05, + 1.883624081529e-05, + 2.016136713792e-05, + 2.150198033632e-05, + 2.285562732141e-05,  \
+ 2.421986500849e-05, + 2.559235435911e-05, + 2.697083837120e-05, + 2.835296400008e-05, + 2.973667033075e-05,  \
+ 3.111963033007e-05, + 3.249973506172e-05, + 3.387491560716e-05, + 3.524332314555e-05, + 3.660289876279e-05,  \
+ 3.795185766649e-05, + 3.928847108909e-05, + 4.061119034304e-05, + 4.191839470877e-05, + 4.320883163018e-05,  \
+ 4.448138861335e-05, + 4.573464902933e-05, + 4.696786854765e-05, + 4.818018278456e-05, + 4.937083940604e-05,  \
+ 5.053927416157e-05, + 5.168495881662e-05, + 5.280774530547e-05, + 5.390729747887e-05, + 5.498336722667e-05,  \
+ 5.603611862171e-05, + 5.706552765332e-05, + 5.807163033751e-05, + 5.905479483772e-05, + 6.001521323924e-05,  \
+ 6.095310563978e-05, + 6.186882819748e-05, + 6.276292115217e-05, + 6.363558059093e-05, + 6.448752283177e-05 ]

* Data table for Id-Vg at Vd = 0.56V
.param vg_data_vd0.56=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.56=[ \
+ 4.744090000000e-10, + 6.878620000000e-10, + 9.973240000000e-10, + 1.445900000000e-09, + 2.096200000000e-09,  \
+ 3.038700000000e-09, + 4.404200000000e-09, + 6.382200000000e-09, + 9.245700000000e-09, + 1.338860000000e-08,  \
+ 1.937610000000e-08, + 2.801710000000e-08, + 4.046190000000e-08, + 5.833190000000e-08, + 8.388660000000e-08,  \
+ 1.202220000000e-07, + 1.714820000000e-07, + 2.430520000000e-07, + 3.416430000000e-07, + 4.752100000000e-07,  \
+ 6.525980000000e-07, + 8.829230000000e-07, + 1.174800000000e-06, + 1.535500000000e-06, + 1.970300000000e-06,  \
+ 2.482300000000e-06, + 3.072500000000e-06, + 3.739600000000e-06, + 4.480900000000e-06, + 5.292600000000e-06,  \
+ 6.170000000000e-06, + 7.108300000000e-06, + 8.102300000000e-06, + 9.147000000000e-06, + 1.023780000000e-05,  \
+ 1.137010000000e-05, + 1.253980000000e-05, + 1.374300000000e-05, + 1.497620000000e-05, + 1.623590000000e-05,  \
+ 1.751910000000e-05, + 1.882290000000e-05, + 2.014470000000e-05, + 2.148180000000e-05, + 2.283190000000e-05,  \
+ 2.419280000000e-05, + 2.556220000000e-05, + 2.693810000000e-05, + 2.831850000000e-05, + 2.970140000000e-05,  \
+ 3.108510000000e-05, + 3.246780000000e-05, + 3.384770000000e-05, + 3.522310000000e-05, + 3.659240000000e-05,  \
+ 3.795410000000e-05, + 3.930650000000e-05, + 4.064820000000e-05, + 4.197780000000e-05, + 4.329380000000e-05,  \
+ 4.459480000000e-05, + 4.587950000000e-05, + 4.714670000000e-05, + 4.839500000000e-05, + 4.962340000000e-05,  \
+ 5.083070000000e-05, + 5.201580000000e-05, + 5.317760000000e-05, + 5.431530000000e-05, + 5.542780000000e-05,  \
+ 5.651450000000e-05, + 5.757440000000e-05, + 5.860690000000e-05, + 5.961130000000e-05, + 6.058700000000e-05,  \
+ 6.153370000000e-05, + 6.245070000000e-05, + 6.333780000000e-05, + 6.419460000000e-05, + 6.502100000000e-05 ]

.param id_pred_data_vd0.56=[ \
+ 4.778605822153e-10, + 6.832605503604e-10, + 9.923688004676e-10, + 1.449163384848e-09, + 2.112682864208e-09,  \
+ 3.065644378353e-09, + 4.429760522839e-09, + 6.388182001160e-09, + 9.214979570515e-09, + 1.331172782670e-08,  \
+ 1.925397242530e-08, + 2.785367115621e-08, + 4.024983695672e-08, + 5.803875296806e-08, + 8.345402306986e-08,  \
+ 1.195874085624e-07, + 1.706208399810e-07, + 2.420092459943e-07, + 3.405396500966e-07, + 4.741909333461e-07,  \
+ 6.517495785374e-07, + 8.822082781990e-07, + 1.174040189653e-06, + 1.534475068183e-06, + 1.968948854483e-06,  \
+ 2.480763832864e-06, + 3.071050814469e-06, + 3.738928426174e-06, + 4.481860014494e-06, + 5.296062372508e-06,  \
+ 6.176908864290e-06, + 7.119314977899e-06, + 8.118061741698e-06, + 9.167974494630e-06, + 1.026415920933e-05,  \
+ 1.140198364737e-05, + 1.257720621652e-05, + 1.378590619424e-05, + 1.502457642346e-05, + 1.628987272852e-05,  \
+ 1.757879828801e-05, + 1.888854778372e-05, + 2.021646563662e-05, + 2.156000322429e-05, + 2.291673619766e-05,  \
+ 2.428429521387e-05, + 2.566036186181e-05, + 2.704263810301e-05, + 2.842893183697e-05, + 2.981702855323e-05,  \
+ 3.120479726931e-05, + 3.259007848101e-05, + 3.397073305678e-05, + 3.534489893354e-05, + 3.671063459478e-05,  \
+ 3.806606575381e-05, + 3.940933442209e-05, + 4.073911230080e-05, + 4.205356177408e-05, + 4.335150937550e-05,  \
+ 4.463154939003e-05, + 4.589254094753e-05, + 4.713365691714e-05, + 4.835380124860e-05, + 4.955238720868e-05,  \
+ 5.072864878457e-05, + 5.188228853513e-05, + 5.301280121785e-05, + 5.411997495685e-05, + 5.520355713088e-05,  \
+ 5.626369034871e-05, + 5.730028089602e-05, + 5.831358139403e-05, + 5.930361221544e-05, + 6.027066672686e-05,  \
+ 6.121523794718e-05, + 6.213738699444e-05, + 6.303782691248e-05, + 6.391668401193e-05, + 6.477467541117e-05 ]

* Data table for Id-Vg at Vd = 0.57V
.param vg_data_vd0.57=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.57=[ \
+ 4.789500000000e-10, + 6.943570000000e-10, + 1.006600000000e-09, + 1.459200000000e-09, + 2.115200000000e-09,  \
+ 3.065800000000e-09, + 4.442900000000e-09, + 6.437400000000e-09, + 9.324500000000e-09, + 1.350080000000e-08,  \
+ 1.953580000000e-08, + 2.824390000000e-08, + 4.078330000000e-08, + 5.878590000000e-08, + 8.452510000000e-08,  \
+ 1.211140000000e-07, + 1.727200000000e-07, + 2.447510000000e-07, + 3.439470000000e-07, + 4.782830000000e-07,  \
+ 6.566210000000e-07, + 8.880880000000e-07, + 1.181300000000e-06, + 1.543400000000e-06, + 1.979900000000e-06,  \
+ 2.493700000000e-06, + 3.085700000000e-06, + 3.754700000000e-06, + 4.498000000000e-06, + 5.311700000000e-06,  \
+ 6.191100000000e-06, + 7.131400000000e-06, + 8.127400000000e-06, + 9.174200000000e-06, + 1.026710000000e-05,  \
+ 1.140150000000e-05, + 1.257330000000e-05, + 1.377870000000e-05, + 1.501400000000e-05, + 1.627600000000e-05,  \
+ 1.756150000000e-05, + 1.886770000000e-05, + 2.019200000000e-05, + 2.153170000000e-05, + 2.288450000000e-05,  \
+ 2.424810000000e-05, + 2.562040000000e-05, + 2.699940000000e-05, + 2.838290000000e-05, + 2.976930000000e-05,  \
+ 3.115650000000e-05, + 3.254290000000e-05, + 3.392660000000e-05, + 3.530620000000e-05, + 3.667980000000e-05,  \
+ 3.804600000000e-05, + 3.940320000000e-05, + 4.074990000000e-05, + 4.208470000000e-05, + 4.340620000000e-05,  \
+ 4.471290000000e-05, + 4.600370000000e-05, + 4.727710000000e-05, + 4.853200000000e-05, + 4.976710000000e-05,  \
+ 5.098140000000e-05, + 5.217380000000e-05, + 5.334310000000e-05, + 5.448850000000e-05, + 5.560900000000e-05,  \
+ 5.670380000000e-05, + 5.777200000000e-05, + 5.881300000000e-05, + 5.982600000000e-05, + 6.081050000000e-05,  \
+ 6.176590000000e-05, + 6.269180000000e-05, + 6.358780000000e-05, + 6.445350000000e-05, + 6.528880000000e-05 ]

.param id_pred_data_vd0.57=[ \
+ 4.824825555749e-10, + 6.897126503258e-10, + 1.001682563562e-09, + 1.462853558287e-09, + 2.132868894833e-09,  \
+ 3.095172145251e-09, + 4.472307750802e-09, + 6.448579776830e-09, + 9.299709482491e-09, + 1.342971851059e-08,  \
+ 1.941796515581e-08, + 2.808239518259e-08, + 4.057021683934e-08, + 5.848945498599e-08, + 8.408878031219e-08,  \
+ 1.204787254494e-07, + 1.718630323921e-07, + 2.437197929339e-07, + 3.428606083844e-07, + 4.772857744229e-07,  \
+ 6.558012637470e-07, + 8.874107584234e-07, + 1.180595413643e-06, + 1.542586558116e-06, + 1.978813390906e-06,  \
+ 2.492567568879e-06, + 3.084962900175e-06, + 3.755106549761e-06, + 4.500437562456e-06, + 5.317127206581e-06,  \
+ 6.200542693477e-06, + 7.145559520723e-06, + 8.146931359079e-06, + 9.199480828102e-06, + 1.029825398291e-05,  \
+ 1.143863695688e-05, + 1.261640987650e-05, + 1.382761103741e-05, + 1.506873493781e-05, + 1.633650417716e-05,  \
+ 1.762792544469e-05, + 1.894023353088e-05, + 2.027076068771e-05, + 2.161706208426e-05, + 2.297674887814e-05,  \
+ 2.434737831209e-05, + 2.572682282334e-05, + 2.711273089517e-05, + 2.850291897630e-05, + 2.989525328303e-05,  \
+ 3.128752745397e-05, + 3.267766576755e-05, + 3.406362360693e-05, + 3.544337501808e-05, + 3.681501846586e-05,  \
+ 3.817667522526e-05, + 3.952659513743e-05, + 4.086313587322e-05, + 4.218476293318e-05, + 4.349003720563e-05,  \
+ 4.477762740862e-05, + 4.604638888850e-05, + 4.729523090646e-05, + 4.852330741414e-05, + 4.972979309969e-05,  \
+ 5.091405342682e-05, + 5.207553680521e-05, + 5.321380776877e-05, + 5.432870457298e-05, + 5.542000326386e-05,  \
+ 5.648757942254e-05, + 5.753148281656e-05, + 5.855182957021e-05, + 5.954886022664e-05, + 6.052268261556e-05,  \
+ 6.147372390842e-05, + 6.240232418349e-05, + 6.330889817036e-05, + 6.419386059861e-05, + 6.505780453153e-05 ]

* Data table for Id-Vg at Vd = 0.58V
.param vg_data_vd0.58=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.58=[ \
+ 4.835250000000e-10, + 7.008990000000e-10, + 1.016000000000e-09, + 1.472600000000e-09, + 2.134300000000e-09,  \
+ 3.093100000000e-09, + 4.481900000000e-09, + 6.493000000000e-09, + 9.403800000000e-09, + 1.361370000000e-08,  \
+ 1.969640000000e-08, + 2.847210000000e-08, + 4.110650000000e-08, + 5.924230000000e-08, + 8.516680000000e-08,  \
+ 1.220110000000e-07, + 1.739640000000e-07, + 2.464580000000e-07, + 3.462580000000e-07, + 4.813650000000e-07,  \
+ 6.606560000000e-07, + 8.932640000000e-07, + 1.187800000000e-06, + 1.551400000000e-06, + 1.989500000000e-06,  \
+ 2.505100000000e-06, + 3.098900000000e-06, + 3.769800000000e-06, + 4.515100000000e-06, + 5.330700000000e-06,  \
+ 6.212100000000e-06, + 7.154400000000e-06, + 8.152400000000e-06, + 9.201300000000e-06, + 1.029610000000e-05,  \
+ 1.143260000000e-05, + 1.260650000000e-05, + 1.381400000000e-05, + 1.505150000000e-05, + 1.631570000000e-05,  \
+ 1.760350000000e-05, + 1.891200000000e-05, + 2.023870000000e-05, + 2.158090000000e-05, + 2.293630000000e-05,  \
+ 2.430260000000e-05, + 2.567780000000e-05, + 2.705960000000e-05, + 2.844630000000e-05, + 2.983580000000e-05,  \
+ 3.122650000000e-05, + 3.261640000000e-05, + 3.400390000000e-05, + 3.538730000000e-05, + 3.676510000000e-05,  \
+ 3.813560000000e-05, + 3.949730000000e-05, + 4.084880000000e-05, + 4.218860000000e-05, + 4.351530000000e-05,  \
+ 4.482750000000e-05, + 4.612400000000e-05, + 4.740330000000e-05, + 4.866440000000e-05, + 4.990600000000e-05,  \
+ 5.112690000000e-05, + 5.232620000000e-05, + 5.350270000000e-05, + 5.465540000000e-05, + 5.578350000000e-05,  \
+ 5.688600000000e-05, + 5.796210000000e-05, + 5.901110000000e-05, + 6.003240000000e-05, + 6.102520000000e-05,  \
+ 6.198900000000e-05, + 6.292340000000e-05, + 6.382790000000e-05, + 6.470220000000e-05, + 6.554600000000e-05 ]

.param id_pred_data_vd0.58=[ \
+ 4.871414427399e-10, + 6.961959408969e-10, + 1.011015449137e-09, + 1.476550872681e-09, + 2.153061635646e-09,  \
+ 3.124713554570e-09, + 4.514941576161e-09, + 6.509221179840e-09, + 9.384888102204e-09, + 1.354853942814e-08,  \
+ 1.958337939811e-08, + 2.831324607655e-08, + 4.089397307894e-08, + 5.894530133332e-08, + 8.473136887233e-08,  \
+ 1.213816929635e-07, + 1.731217071210e-07, + 2.454534734397e-07, + 3.452119403846e-07, + 4.804192190022e-07,  \
+ 6.598977142858e-07, + 8.926644977691e-07, + 1.187205507449e-06, + 1.550753127049e-06, + 1.988724061448e-06,  \
+ 2.504413514544e-06, + 3.098905908701e-06, + 3.771301580855e-06, + 4.519002031884e-06, + 5.338169648894e-06,  \
+ 6.224125972949e-06, + 7.171738361649e-06, + 8.175710645446e-06, + 9.230860596290e-06, + 1.033218850353e-05,  \
+ 1.147511455201e-05, + 1.265533956030e-05, + 1.386898213241e-05, + 1.511249320174e-05, + 1.638266236114e-05,  \
+ 1.767648598616e-05, + 1.899119466543e-05, + 2.032425531070e-05, + 2.167313694372e-05, + 2.303551642399e-05,  \
+ 2.440911703161e-05, + 2.579164305644e-05, + 2.718096548051e-05, + 2.857478648366e-05, + 2.997108887939e-05,  \
+ 3.136764236842e-05, + 3.276246563473e-05, + 3.415338956984e-05, + 3.553853413905e-05, + 3.691587160574e-05,  \
+ 3.828359156614e-05, + 3.963990049670e-05, + 4.098312725546e-05, + 4.231174418237e-05, + 4.362427425804e-05,  \
+ 4.491930798395e-05, + 4.619569750503e-05, + 4.745238780743e-05, + 4.868830699706e-05, + 4.990270390408e-05,  \
+ 5.109492863994e-05, + 5.226432709605e-05, + 5.341059542843e-05, + 5.453330741148e-05, + 5.563227314269e-05,  \
+ 5.670745464158e-05, + 5.775872108643e-05, + 5.878635100089e-05, + 5.979034016491e-05, + 6.077106838347e-05,  \
+ 6.172871711897e-05, + 6.266374213737e-05, + 6.357654012390e-05, + 6.446751620388e-05, + 6.533726540511e-05 ]

* Data table for Id-Vg at Vd = 0.59V
.param vg_data_vd0.59=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.59=[ \
+ 4.881350000000e-10, + 7.074910000000e-10, + 1.025400000000e-09, + 1.486100000000e-09, + 2.153500000000e-09,  \
+ 3.120500000000e-09, + 4.521100000000e-09, + 6.548900000000e-09, + 9.483500000000e-09, + 1.372730000000e-08,  \
+ 1.985800000000e-08, + 2.870150000000e-08, + 4.143140000000e-08, + 5.970120000000e-08, + 8.581180000000e-08,  \
+ 1.229120000000e-07, + 1.752130000000e-07, + 2.481720000000e-07, + 3.485780000000e-07, + 4.844560000000e-07,  \
+ 6.647010000000e-07, + 8.984510000000e-07, + 1.194300000000e-06, + 1.559400000000e-06, + 1.999200000000e-06,  \
+ 2.516500000000e-06, + 3.112100000000e-06, + 3.784900000000e-06, + 4.532100000000e-06, + 5.349700000000e-06,  \
+ 6.233100000000e-06, + 7.177300000000e-06, + 8.177300000000e-06, + 9.228200000000e-06, + 1.032510000000e-05,  \
+ 1.146360000000e-05, + 1.263950000000e-05, + 1.384910000000e-05, + 1.508870000000e-05, + 1.635510000000e-05,  \
+ 1.764510000000e-05, + 1.895590000000e-05, + 2.028490000000e-05, + 2.162950000000e-05, + 2.298750000000e-05,  \
+ 2.435640000000e-05, + 2.573430000000e-05, + 2.711900000000e-05, + 2.850860000000e-05, + 2.990120000000e-05,  \
+ 3.129510000000e-05, + 3.268840000000e-05, + 3.407950000000e-05, + 3.546670000000e-05, + 3.684840000000e-05,  \
+ 3.822300000000e-05, + 3.958910000000e-05, + 4.094510000000e-05, + 4.228970000000e-05, + 4.362130000000e-05,  \
+ 4.493870000000e-05, + 4.624060000000e-05, + 4.752560000000e-05, + 4.879260000000e-05, + 5.004030000000e-05,  \
+ 5.126760000000e-05, + 5.247340000000e-05, + 5.365660000000e-05, + 5.481630000000e-05, + 5.595160000000e-05,  \
+ 5.706140000000e-05, + 5.814510000000e-05, + 5.920180000000e-05, + 6.023090000000e-05, + 6.123160000000e-05,  \
+ 6.220350000000e-05, + 6.314600000000e-05, + 6.405860000000e-05, + 6.494110000000e-05, + 6.579300000000e-05 ]

.param id_pred_data_vd0.59=[ \
+ 4.918379326035e-10, + 7.027135606741e-10, + 1.020365428817e-09, + 1.490248864311e-09, + 2.173242961145e-09,  \
+ 3.154261101201e-09, + 4.557643737968e-09, + 6.570033344033e-09, + 9.470488571139e-09, + 1.366807559577e-08,  \
+ 1.975001975296e-08, + 2.854600186453e-08, + 4.122071210588e-08, + 5.940585197095e-08, + 8.538125626956e-08,  \
+ 1.222956503000e-07, + 1.743961456668e-07, + 2.472092134553e-07, + 3.475927178442e-07, + 4.835890632648e-07,  \
+ 6.640383128342e-07, + 8.979683570942e-07, + 1.193866594349e-06, + 1.558966216635e-06, + 1.998683012516e-06,  \
+ 2.516292265682e-06, + 3.112871204394e-06, + 3.787491373259e-06, + 4.537545155472e-06, + 5.359169017538e-06,  \
+ 6.247644887480e-06, + 7.197815484687e-06, + 8.204358255171e-06, + 9.262066014344e-06, + 1.036592153469e-05,  \
+ 1.151132721134e-05, + 1.269398057048e-05, + 1.391001593220e-05, + 1.515584772278e-05, + 1.642828208787e-05,  \
+ 1.772440635250e-05, + 1.904142482090e-05, + 2.037678863417e-05, + 2.172810025513e-05, + 2.309305444214e-05,  \
+ 2.446933951433e-05, + 2.585480691778e-05, + 2.724724370637e-05, + 2.864454640076e-05, + 3.004454498296e-05,  \
+ 3.144518319459e-05, + 3.284432965302e-05, + 3.423996888159e-05, + 3.563022492017e-05, + 3.701302004629e-05,  \
+ 3.838657059532e-05, + 3.974907143856e-05, + 4.109877969313e-05, + 4.243421863066e-05, + 4.375376127427e-05,  \
+ 4.505616270762e-05, + 4.634010932932e-05, + 4.760445066495e-05, + 4.884828951617e-05, + 5.007068575651e-05,  \
+ 5.127093536430e-05, + 5.244836436759e-05, + 5.360265509808e-05, + 5.473326666106e-05, + 5.584015183558e-05,  \
+ 5.692303588148e-05, + 5.798189733468e-05, + 5.901681775867e-05, + 6.002800750139e-05, + 6.101565544668e-05,  \
+ 6.198011789820e-05, + 6.292164813203e-05, + 6.384064108715e-05, + 6.473772780737e-05, + 6.561324742506e-05 ]

* Data table for Id-Vg at Vd = 0.60V
.param vg_data_vd0.60=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.60=[ \
+ 4.927800000000e-10, + 7.141320000000e-10, + 1.034900000000e-09, + 1.499600000000e-09, + 2.172900000000e-09,  \
+ 3.148200000000e-09, + 4.560600000000e-09, + 6.605200000000e-09, + 9.563800000000e-09, + 1.384160000000e-08,  \
+ 2.002050000000e-08, + 2.893220000000e-08, + 4.175820000000e-08, + 6.016250000000e-08, + 8.646010000000e-08,  \
+ 1.238180000000e-07, + 1.764680000000e-07, + 2.498920000000e-07, + 3.509070000000e-07, + 4.875590000000e-07,  \
+ 6.687580000000e-07, + 9.036500000000e-07, + 1.200800000000e-06, + 1.567400000000e-06, + 2.008800000000e-06,  \
+ 2.527800000000e-06, + 3.125300000000e-06, + 3.800000000000e-06, + 4.549100000000e-06, + 5.368600000000e-06,  \
+ 6.254000000000e-06, + 7.200200000000e-06, + 8.202200000000e-06, + 9.255000000000e-06, + 1.035380000000e-05,  \
+ 1.149430000000e-05, + 1.267230000000e-05, + 1.388390000000e-05, + 1.512560000000e-05, + 1.639410000000e-05,  \
+ 1.768630000000e-05, + 1.899930000000e-05, + 2.033060000000e-05, + 2.167760000000e-05, + 2.303800000000e-05,  \
+ 2.440950000000e-05, + 2.578990000000e-05, + 2.717740000000e-05, + 2.856990000000e-05, + 2.996550000000e-05,  \
+ 3.136250000000e-05, + 3.275910000000e-05, + 3.415360000000e-05, + 3.554440000000e-05, + 3.692980000000e-05,  \
+ 3.830840000000e-05, + 3.967860000000e-05, + 4.103900000000e-05, + 4.238810000000e-05, + 4.372450000000e-05,  \
+ 4.504690000000e-05, + 4.635390000000e-05, + 4.764430000000e-05, + 4.891680000000e-05, + 5.017030000000e-05,  \
+ 5.140370000000e-05, + 5.261570000000e-05, + 5.380540000000e-05, + 5.497170000000e-05, + 5.611380000000e-05,  \
+ 5.723070000000e-05, + 5.832150000000e-05, + 5.938550000000e-05, + 6.042200000000e-05, + 6.143040000000e-05,  \
+ 6.240990000000e-05, + 6.336010000000e-05, + 6.428060000000e-05, + 6.517090000000e-05, + 6.603070000000e-05 ]

.param id_pred_data_vd0.60=[ \
+ 4.965734157203e-10, + 7.092601839176e-10, + 1.029731899749e-09, + 1.503940172398e-09, + 2.193393067174e-09,  \
+ 3.183768448878e-09, + 4.600340908212e-09, + 6.630962978704e-09, + 9.556348246065e-09, + 1.378820257969e-08,  \
+ 1.991767177856e-08, + 2.878063654066e-08, + 4.155033224151e-08, + 5.987083682157e-08, + 8.603798846707e-08,  \
+ 1.232199792867e-07, + 1.756859489888e-07, + 2.489859923571e-07, + 3.500015168356e-07, + 4.867945108344e-07,  \
+ 6.682199455099e-07, + 9.033164360517e-07, + 1.200573797178e-06, + 1.567222443555e-06, + 2.008672072407e-06,  \
+ 2.528188269935e-06, + 3.126826959488e-06, + 3.803659092227e-06, + 4.556041039905e-06, + 5.380085531215e-06,  \
+ 6.271054007811e-06, + 7.223744069051e-06, + 8.232837899413e-06, + 9.293064067606e-06, + 1.039942399075e-05,  \
+ 1.154725359811e-05, + 1.273227571801e-05, + 1.395059516653e-05, + 1.519868455944e-05, + 1.647333192523e-05,  \
+ 1.777162106009e-05, + 1.909080165206e-05, + 2.042836131295e-05, + 2.178195136366e-05, + 2.314927114639e-05,  \
+ 2.452806365909e-05, + 2.591621378087e-05, + 2.731159547693e-05, + 2.871203250834e-05, + 3.011544467881e-05,  \
+ 3.151986747980e-05, + 3.292312248959e-05, + 3.432325611357e-05, + 3.571829074644e-05, + 3.710630990099e-05,  \
+ 3.848537744489e-05, + 3.985385410488e-05, + 4.120987141505e-05, + 4.255188396201e-05, + 4.387843364384e-05,  \
+ 4.518794885371e-05, + 4.647937312257e-05, + 4.775138804689e-05, + 4.900298954453e-05, + 5.023337871535e-05,  \
+ 5.144164751982e-05, + 5.262721097097e-05, + 5.378959758673e-05, + 5.492828786373e-05, + 5.604306788882e-05,  \
+ 5.713381542591e-05, + 5.820036894875e-05, + 5.924297729507e-05, + 6.026148766978e-05, + 6.125619256636e-05,  \
+ 6.222754163900e-05, + 6.317578372546e-05, + 6.410123314708e-05, + 6.500440067612e-05, + 6.588591495529e-05 ]

* Data table for Id-Vg at Vd = 0.61V
.param vg_data_vd0.61=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.61=[ \
+ 4.974610000000e-10, + 7.208220000000e-10, + 1.044400000000e-09, + 1.513300000000e-09, + 2.192400000000e-09,  \
+ 3.176000000000e-09, + 4.600300000000e-09, + 6.661900000000e-09, + 9.644600000000e-09, + 1.395660000000e-08,  \
+ 2.018400000000e-08, + 2.916430000000e-08, + 4.208690000000e-08, + 6.062630000000e-08, + 8.711180000000e-08,  \
+ 1.247280000000e-07, + 1.777290000000e-07, + 2.516200000000e-07, + 3.532450000000e-07, + 4.906710000000e-07,  \
+ 6.728270000000e-07, + 9.088610000000e-07, + 1.207300000000e-06, + 1.575500000000e-06, + 2.018400000000e-06,  \
+ 2.539200000000e-06, + 3.138500000000e-06, + 3.815100000000e-06, + 4.566000000000e-06, + 5.387500000000e-06,  \
+ 6.274800000000e-06, + 7.222900000000e-06, + 8.226900000000e-06, + 9.281600000000e-06, + 1.038250000000e-05,  \
+ 1.152500000000e-05, + 1.270490000000e-05, + 1.391850000000e-05, + 1.516230000000e-05, + 1.643280000000e-05,  \
+ 1.772710000000e-05, + 1.904230000000e-05, + 2.037590000000e-05, + 2.172520000000e-05, + 2.308790000000e-05,  \
+ 2.446180000000e-05, + 2.584490000000e-05, + 2.723500000000e-05, + 2.863020000000e-05, + 3.002870000000e-05,  \
+ 3.142870000000e-05, + 3.282850000000e-05, + 3.422630000000e-05, + 3.562050000000e-05, + 3.700960000000e-05,  \
+ 3.839200000000e-05, + 3.976610000000e-05, + 4.113060000000e-05, + 4.248400000000e-05, + 4.382490000000e-05,  \
+ 4.515200000000e-05, + 4.646400000000e-05, + 4.775950000000e-05, + 4.903740000000e-05, + 5.029640000000e-05,  \
+ 5.153550000000e-05, + 5.275350000000e-05, + 5.394930000000e-05, + 5.512200000000e-05, + 5.627050000000e-05,  \
+ 5.739400000000e-05, + 5.849170000000e-05, + 5.956270000000e-05, + 6.060640000000e-05, + 6.162190000000e-05,  \
+ 6.260880000000e-05, + 6.356640000000e-05, + 6.449430000000e-05, + 6.539210000000e-05, + 6.625940000000e-05 ]

.param id_pred_data_vd0.61=[ \
+ 5.013510040452e-10, + 7.158382286931e-10, + 1.039109743806e-09, + 1.517610532797e-09, + 2.213490886138e-09,  \
+ 3.213216577258e-09, + 4.642998128190e-09, + 6.691913476686e-09, + 9.642403373533e-09, + 1.390881058327e-08,  \
+ 2.008626413641e-08, + 2.901671905420e-08, + 4.188245718240e-08, + 6.033996321264e-08, + 8.670122781496e-08,  \
+ 1.241538677732e-07, + 1.769899645865e-07, + 2.507828870080e-07, + 3.524363251017e-07, + 4.900332481839e-07,  \
+ 6.724406330250e-07, + 9.087073760838e-07, + 1.207321895436e-06, + 1.575515832428e-06, + 2.018687241616e-06,  \
+ 2.540088867136e-06, + 3.140778558191e-06, + 3.819785429187e-06, + 4.574458407660e-06, + 5.400891204772e-06,  \
+ 6.294315107880e-06, + 7.249508971654e-06, + 8.261082439276e-06, + 9.323799386038e-06, + 1.043260399456e-05,  \
+ 1.158282602773e-05, + 1.277015808228e-05, + 1.399072882123e-05, + 1.524099867311e-05, + 1.651774540733e-05,  \
+ 1.781807301086e-05, + 1.913929740113e-05, + 2.047894420684e-05, + 2.183461561799e-05, + 2.320411465917e-05,  \
+ 2.458521328663e-05, + 2.597582770250e-05, + 2.737381862971e-05, + 2.877717328374e-05, + 3.018382562004e-05,  \
+ 3.159167852573e-05, + 3.299873031210e-05, + 3.440309468715e-05, + 3.580263681215e-05, + 3.719556360011e-05,  \
+ 3.857997544401e-05, + 3.995406150352e-05, + 4.131608860916e-05, + 4.266452997399e-05, + 4.399777892104e-05,  \
+ 4.531435748504e-05, + 4.661304068577e-05, + 4.789268787135e-05, + 4.915206962323e-05, + 5.039028495958e-05,  \
+ 5.160661043192e-05, + 5.280035809847e-05, + 5.397084001743e-05, + 5.511767893040e-05, + 5.624064848234e-05,  \
+ 5.733939360653e-05, + 5.841385216627e-05, + 5.946408185991e-05, + 6.049020252249e-05, + 6.149237837235e-05,  \
+ 6.247074699786e-05, + 6.342572116409e-05, + 6.435784234782e-05, + 6.526742567075e-05, + 6.615490165132e-05 ]

* Data table for Id-Vg at Vd = 0.62V
.param vg_data_vd0.62=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.62=[ \
+ 5.021770000000e-10, + 7.275630000000e-10, + 1.054100000000e-09, + 1.527000000000e-09, + 2.212100000000e-09,  \
+ 3.204100000000e-09, + 4.640300000000e-09, + 6.719000000000e-09, + 9.725900000000e-09, + 1.407230000000e-08,  \
+ 2.034850000000e-08, + 2.939780000000e-08, + 4.241740000000e-08, + 6.109270000000e-08, + 8.776680000000e-08,  \
+ 1.256420000000e-07, + 1.789950000000e-07, + 2.533560000000e-07, + 3.555910000000e-07, + 4.937940000000e-07,  \
+ 6.769070000000e-07, + 9.140850000000e-07, + 1.213900000000e-06, + 1.583500000000e-06, + 2.028100000000e-06,  \
+ 2.550600000000e-06, + 3.151700000000e-06, + 3.830100000000e-06, + 4.583000000000e-06, + 5.406400000000e-06,  \
+ 6.295600000000e-06, + 7.245700000000e-06, + 8.251500000000e-06, + 9.308200000000e-06, + 1.041100000000e-05,  \
+ 1.155540000000e-05, + 1.273730000000e-05, + 1.395290000000e-05, + 1.519860000000e-05, + 1.647120000000e-05,  \
+ 1.776760000000e-05, + 1.908500000000e-05, + 2.042070000000e-05, + 2.177220000000e-05, + 2.313720000000e-05,  \
+ 2.451360000000e-05, + 2.589910000000e-05, + 2.729180000000e-05, + 2.868970000000e-05, + 3.009100000000e-05,  \
+ 3.149390000000e-05, + 3.289670000000e-05, + 3.429760000000e-05, + 3.569520000000e-05, + 3.708770000000e-05,  \
+ 3.847370000000e-05, + 3.985170000000e-05, + 4.122010000000e-05, + 4.257770000000e-05, + 4.392290000000e-05,  \
+ 4.525450000000e-05, + 4.657110000000e-05, + 4.787160000000e-05, + 4.915450000000e-05, + 5.041880000000e-05,  \
+ 5.166340000000e-05, + 5.288700000000e-05, + 5.408860000000e-05, + 5.526730000000e-05, + 5.642210000000e-05,  \
+ 5.755200000000e-05, + 5.865610000000e-05, + 5.973380000000e-05, + 6.078420000000e-05, + 6.180670000000e-05,  \
+ 6.280050000000e-05, + 6.376520000000e-05, + 6.470030000000e-05, + 6.560520000000e-05, + 6.647970000000e-05 ]

.param id_pred_data_vd0.62=[ \
+ 5.061688279628e-10, + 7.224484654955e-10, + 1.048497166867e-09, + 1.531256539344e-09, + 2.233530360662e-09,  \
+ 3.242573010098e-09, + 4.685568750773e-09, + 6.752845180813e-09, + 9.728549166255e-09, + 1.402975367881e-08,  \
+ 2.025555090768e-08, + 2.925407272869e-08, + 4.221675780514e-08, + 6.081265794933e-08, + 8.736993805769e-08,  \
+ 1.250965320310e-07, + 1.783067415317e-07, + 2.525978470658e-07, + 3.548952497567e-07, + 4.933015611641e-07,  \
+ 6.766970454919e-07, + 9.141332475338e-07, + 1.214104627252e-06, + 1.583835278325e-06, + 2.028716098721e-06,  \
+ 2.551987463448e-06, + 3.154693549732e-06, + 3.835848965537e-06, + 4.592784553097e-06, + 5.421566638688e-06,  \
+ 6.317398238025e-06, + 7.275040279637e-06, + 8.289092984342e-06, + 9.354236080981e-06, + 1.046543293342e-05,  \
+ 1.161798805697e-05, + 1.280759392102e-05, + 1.403033715178e-05, + 1.528265962406e-05, + 1.656144417211e-05,  \
+ 1.786372926290e-05, + 1.918689282320e-05, + 2.052842442936e-05, + 2.188603357354e-05, + 2.325755944184e-05,  \
+ 2.464073520969e-05, + 2.603357148473e-05, + 2.743401571934e-05, + 2.883998829930e-05, + 3.024951111001e-05,  \
+ 3.166057897033e-05, + 3.307120248792e-05, + 3.447937648161e-05, + 3.588311607018e-05, + 3.728063260496e-05,  \
+ 3.867005172651e-05, + 4.004952614196e-05, + 4.141741155763e-05, + 4.277193511371e-05, + 4.411173897097e-05,  \
+ 4.543514951365e-05, + 4.674099385738e-05, + 4.802799987374e-05, + 4.929507587804e-05, + 5.054113920778e-05,  \
+ 5.176549966563e-05, + 5.296726405504e-05, + 5.414599028882e-05, + 5.530113703571e-05, + 5.643225769745e-05,  \
+ 5.753913574154e-05, + 5.862175763468e-05, + 5.967987977783e-05, + 6.071377283661e-05, + 6.172347741085e-05,  \
+ 6.270923709963e-05, + 6.367137670168e-05, + 6.461024808232e-05, + 6.552633392857e-05, + 6.642012143857e-05 ]

* Data table for Id-Vg at Vd = 0.63V
.param vg_data_vd0.63=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.63=[ \
+ 5.069300000000e-10, + 7.343550000000e-10, + 1.063800000000e-09, + 1.540900000000e-09, + 2.231900000000e-09,  \
+ 3.232300000000e-09, + 4.680600000000e-09, + 6.776400000000e-09, + 9.807700000000e-09, + 1.418870000000e-08,  \
+ 2.051410000000e-08, + 2.963260000000e-08, + 4.274980000000e-08, + 6.156150000000e-08, + 8.842520000000e-08,  \
+ 1.265610000000e-07, + 1.802670000000e-07, + 2.550980000000e-07, + 3.579470000000e-07, + 4.969280000000e-07,  \
+ 6.809990000000e-07, + 9.193200000000e-07, + 1.220400000000e-06, + 1.591500000000e-06, + 2.037700000000e-06,  \
+ 2.562000000000e-06, + 3.164900000000e-06, + 3.845100000000e-06, + 4.599900000000e-06, + 5.425200000000e-06,  \
+ 6.316300000000e-06, + 7.268300000000e-06, + 8.276100000000e-06, + 9.334600000000e-06, + 1.043930000000e-05,  \
+ 1.158570000000e-05, + 1.276950000000e-05, + 1.398710000000e-05, + 1.523480000000e-05, + 1.650940000000e-05,  \
+ 1.780780000000e-05, + 1.912720000000e-05, + 2.046500000000e-05, + 2.181880000000e-05, + 2.318600000000e-05,  \
+ 2.456470000000e-05, + 2.595260000000e-05, + 2.734780000000e-05, + 2.874830000000e-05, + 3.015230000000e-05,  \
+ 3.155800000000e-05, + 3.296370000000e-05, + 3.436770000000e-05, + 3.576850000000e-05, + 3.716430000000e-05,  \
+ 3.855380000000e-05, + 3.993540000000e-05, + 4.130760000000e-05, + 4.266910000000e-05, + 4.401850000000e-05,  \
+ 4.535440000000e-05, + 4.667550000000e-05, + 4.798060000000e-05, + 4.926840000000e-05, + 5.053780000000e-05,  \
+ 5.178750000000e-05, + 5.301650000000e-05, + 5.422370000000e-05, + 5.540810000000e-05, + 5.656880000000e-05,  \
+ 5.770470000000e-05, + 5.881510000000e-05, + 5.989920000000e-05, + 6.095600000000e-05, + 6.198500000000e-05,  \
+ 6.298560000000e-05, + 6.395710000000e-05, + 6.489890000000e-05, + 6.581080000000e-05, + 6.669210000000e-05 ]

.param id_pred_data_vd0.63=[ \
+ 5.110306078304e-10, + 7.290913972557e-10, + 1.057891874101e-09, + 1.544870751324e-09, + 2.253491553361e-09,  \
+ 3.271813979744e-09, + 4.728011901989e-09, + 6.813663473437e-09, + 9.814745016712e-09, + 1.415087327317e-08,  \
+ 2.042527651014e-08, + 2.949239124916e-08, + 4.255288153843e-08, + 6.128842393593e-08, + 8.804406675722e-08,  \
+ 1.260474425635e-07, + 1.796359285322e-07, + 2.544296242490e-07, + 3.573768276510e-07, + 4.965960442860e-07,  \
+ 6.809824742504e-07, + 9.195907318826e-07, + 1.220914052737e-06, + 1.592171647644e-06, + 2.038742525201e-06,  \
+ 2.563861453382e-06, + 3.168553066644e-06, + 3.851822812067e-06, + 4.610977962329e-06, + 5.442072679216e-06,  \
+ 6.340270711007e-06, + 7.300307788682e-06, + 8.316772100443e-06, + 9.384317154399e-06, + 1.049786633303e-05,  \
+ 1.165269368357e-05, + 1.284449210289e-05, + 1.406932291502e-05, + 1.532367832624e-05, + 1.660438974795e-05,  \
+ 1.790851549231e-05, + 1.923345422256e-05, + 2.057677076664e-05, + 2.193617663579e-05, + 2.330946470465e-05,  \
+ 2.469454931997e-05, + 2.608940900245e-05, + 2.749201768893e-05, + 2.890041119826e-05, + 3.031254054804e-05,  \
+ 3.172648739564e-05, + 3.314026922453e-05, + 3.455200894678e-05, + 3.595970112656e-05, + 3.736155347724e-05,  \
+ 3.875565453200e-05, + 4.014024409116e-05, + 4.151357112278e-05, + 4.287393501727e-05, + 4.421988269314e-05,  \
+ 4.555001607514e-05, + 4.686278123700e-05, + 4.815699554456e-05, + 4.943153136992e-05, + 5.068543985544e-05,  \
+ 5.191780423047e-05, + 5.312761146342e-05, + 5.431461861008e-05, + 5.547796848987e-05, + 5.661740440701e-05,  \
+ 5.773259174020e-05, + 5.882345256396e-05, + 5.988972559862e-05, + 6.093161711760e-05, + 6.194907669851e-05,  \
+ 6.294240229181e-05, + 6.391195602191e-05, + 6.485790290753e-05, + 6.578088927199e-05, + 6.668107096630e-05 ]

* Data table for Id-Vg at Vd = 0.64V
.param vg_data_vd0.64=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.64=[ \
+ 5.117200000000e-10, + 7.411980000000e-10, + 1.073500000000e-09, + 1.554900000000e-09, + 2.251800000000e-09,  \
+ 3.260800000000e-09, + 4.721200000000e-09, + 6.834200000000e-09, + 9.890000000000e-09, + 1.430590000000e-08,  \
+ 2.068060000000e-08, + 2.986890000000e-08, + 4.308410000000e-08, + 6.203300000000e-08, + 8.908720000000e-08,  \
+ 1.274850000000e-07, + 1.815450000000e-07, + 2.568480000000e-07, + 3.603120000000e-07, + 5.000720000000e-07,  \
+ 6.851030000000e-07, + 9.245690000000e-07, + 1.227000000000e-06, + 1.599600000000e-06, + 2.047400000000e-06,  \
+ 2.573400000000e-06, + 3.178100000000e-06, + 3.860200000000e-06, + 4.616800000000e-06, + 5.444000000000e-06,  \
+ 6.337000000000e-06, + 7.290900000000e-06, + 8.300500000000e-06, + 9.361000000000e-06, + 1.046760000000e-05,  \
+ 1.161580000000e-05, + 1.280160000000e-05, + 1.402100000000e-05, + 1.527070000000e-05, + 1.654720000000e-05,  \
+ 1.784760000000e-05, + 1.916910000000e-05, + 2.050900000000e-05, + 2.186490000000e-05, + 2.323430000000e-05,  \
+ 2.461530000000e-05, + 2.600550000000e-05, + 2.740310000000e-05, + 2.880610000000e-05, + 3.021270000000e-05,  \
+ 3.162110000000e-05, + 3.302970000000e-05, + 3.443660000000e-05, + 3.584040000000e-05, + 3.723950000000e-05,  \
+ 3.863230000000e-05, + 4.001740000000e-05, + 4.139330000000e-05, + 4.275850000000e-05, + 4.411190000000e-05,  \
+ 4.545190000000e-05, + 4.677730000000e-05, + 4.808680000000e-05, + 4.937930000000e-05, + 5.065340000000e-05,  \
+ 5.190810000000e-05, + 5.314230000000e-05, + 5.435480000000e-05, + 5.554470000000e-05, + 5.671100000000e-05,  \
+ 5.785270000000e-05, + 5.896900000000e-05, + 6.005910000000e-05, + 6.112220000000e-05, + 6.215750000000e-05,  \
+ 6.316440000000e-05, + 6.414230000000e-05, + 6.509070000000e-05, + 6.600910000000e-05, + 6.689710000000e-05 ]

.param id_pred_data_vd0.64=[ \
+ 5.159360227935e-10, + 7.357671449881e-10, + 1.067293169399e-09, + 1.558451145911e-09, + 2.273361872085e-09,  \
+ 3.300915238924e-09, + 4.770283794642e-09, + 6.874320206407e-09, + 9.900795703288e-09, + 1.427200118087e-08,  \
+ 2.059531880150e-08, + 2.973145228680e-08, + 4.289044682082e-08, + 6.176683655212e-08, + 8.872236321622e-08,  \
+ 1.270053235203e-07, + 1.809756759030e-07, + 2.562760892033e-07, + 3.598777402658e-07, + 4.999148222851e-07,  \
+ 6.852923252154e-07, + 9.250727453036e-07, + 1.227742613992e-06, + 1.600513351150e-06, + 2.048755559372e-06,  \
+ 2.575691905804e-06, + 3.182339132763e-06, + 3.867681662086e-06, + 4.629017785192e-06, + 5.462353001349e-06,  \
+ 6.362878484651e-06, + 7.325269980356e-06, + 8.344087982550e-06, + 9.413963416591e-06, + 1.052981475368e-05,  \
+ 1.168686314486e-05, + 1.288079423830e-05, + 1.410767319612e-05, + 1.536395284347e-05, + 1.664649113081e-05,  \
+ 1.795238233171e-05, + 1.927902339958e-05, + 2.062392653897e-05, + 2.198494039476e-05, + 2.335990080610e-05,  \
+ 2.474665874615e-05, + 2.614331431687e-05, + 2.754785120487e-05, + 2.895830431953e-05, + 3.037279704586e-05,  \
+ 3.178937360644e-05, + 3.320605261251e-05, + 3.462099004537e-05, + 3.603231860325e-05, + 3.743810812011e-05,  \
+ 3.883654484525e-05, + 4.022583365440e-05, + 4.160438198596e-05, + 4.297039005905e-05, + 4.432236775756e-05,  \
+ 4.565871320665e-05, + 4.697815515101e-05, + 4.827946890146e-05, + 4.956135991961e-05, + 5.082292016596e-05,  \
+ 5.206304602325e-05, + 5.328101571649e-05, + 5.447617731988e-05, + 5.564792081714e-05, + 5.679566878825e-05,  \
+ 5.791928619146e-05, + 5.901845637709e-05, + 6.009296514094e-05, + 6.114311050624e-05, + 6.216849200428e-05,  \
+ 6.316972896457e-05, + 6.414688657969e-05, + 6.510028615594e-05, + 6.603030953556e-05, + 6.693741772324e-05 ]

* Data table for Id-Vg at Vd = 0.65V
.param vg_data_vd0.65=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.65=[ \
+ 5.165460000000e-10, + 7.480930000000e-10, + 1.083400000000e-09, + 1.568900000000e-09, + 2.271800000000e-09,  \
+ 3.289400000000e-09, + 4.762000000000e-09, + 6.892400000000e-09, + 9.972900000000e-09, + 1.442380000000e-08,  \
+ 2.084810000000e-08, + 3.010650000000e-08, + 4.342030000000e-08, + 6.250710000000e-08, + 8.975260000000e-08,  \
+ 1.284130000000e-07, + 1.828290000000e-07, + 2.586060000000e-07, + 3.626860000000e-07, + 5.032280000000e-07,  \
+ 6.892200000000e-07, + 9.298310000000e-07, + 1.233600000000e-06, + 1.607600000000e-06, + 2.057100000000e-06,  \
+ 2.584700000000e-06, + 3.191200000000e-06, + 3.875200000000e-06, + 4.633700000000e-06, + 5.462700000000e-06,  \
+ 6.357600000000e-06, + 7.313400000000e-06, + 8.324900000000e-06, + 9.387300000000e-06, + 1.049570000000e-05,  \
+ 1.164580000000e-05, + 1.283350000000e-05, + 1.405480000000e-05, + 1.530630000000e-05, + 1.658480000000e-05,  \
+ 1.788720000000e-05, + 1.921070000000e-05, + 2.055260000000e-05, + 2.191050000000e-05, + 2.328220000000e-05,  \
+ 2.466530000000e-05, + 2.605780000000e-05, + 2.745780000000e-05, + 2.886320000000e-05, + 3.027230000000e-05,  \
+ 3.168340000000e-05, + 3.309460000000e-05, + 3.450440000000e-05, + 3.591120000000e-05, + 3.731330000000e-05,  \
+ 3.870930000000e-05, + 4.009780000000e-05, + 4.147710000000e-05, + 4.284610000000e-05, + 4.420320000000e-05,  \
+ 4.554710000000e-05, + 4.687660000000e-05, + 4.819040000000e-05, + 4.948730000000e-05, + 5.076600000000e-05,  \
+ 5.202550000000e-05, + 5.326460000000e-05, + 5.448220000000e-05, + 5.567730000000e-05, + 5.684890000000e-05,  \
+ 5.799620000000e-05, + 5.911820000000e-05, + 6.021400000000e-05, + 6.128300000000e-05, + 6.232430000000e-05,  \
+ 6.333730000000e-05, + 6.432140000000e-05, + 6.527610000000e-05, + 6.620080000000e-05, + 6.709510000000e-05 ]

.param id_pred_data_vd0.65=[ \
+ 5.208905168308e-10, + 7.424784953525e-10, + 1.076697897506e-09, + 1.571988816895e-09, + 2.293136136533e-09,  \
+ 3.329856057555e-09, + 4.812355269834e-09, + 6.934776042300e-09, + 9.986686499985e-09, + 1.439306798190e-08,  \
+ 2.076550824626e-08, + 2.997107930724e-08, + 4.322911983934e-08, + 6.224744133476e-08, + 8.940469413687e-08,  \
+ 1.279693734091e-07, + 1.823239955456e-07, + 2.581359652254e-07, + 3.623951101872e-07, + 5.032528548554e-07,  \
+ 6.896247498389e-07, + 9.305714229413e-07, + 1.234578661524e-06, + 1.608847969692e-06, + 2.058743120870e-06,  \
+ 2.587468338788e-06, + 3.196023294549e-06, + 3.883390877490e-06, + 4.646852880796e-06, + 5.482394954015e-06,  \
+ 6.385189590219e-06, + 7.349868656092e-06, + 8.370982732231e-06, + 9.443144472243e-06, + 1.056122546288e-05,  \
+ 1.172043012048e-05, + 1.291643402510e-05, + 1.414527750967e-05, + 1.540340763313e-05, + 1.668768054515e-05,  \
+ 1.799522315196e-05, + 1.932337163453e-05, + 2.066985234705e-05, + 2.203229705628e-05, + 2.340867922612e-05,  \
+ 2.479701015545e-05, + 2.619523493195e-05, + 2.760145234788e-05, + 2.901373754867e-05, + 3.043032884307e-05,  \
+ 3.184916186001e-05, + 3.326850564918e-05, + 3.468630529824e-05, + 3.610087951529e-05, + 3.751027506951e-05,  \
+ 3.891274445778e-05, + 4.030648342450e-05, + 4.168982959527e-05, + 4.306110640755e-05, + 4.441864912224e-05,  \
+ 4.576108622132e-05, + 4.708711712738e-05, + 4.839514331252e-05, + 4.968417633791e-05, + 5.095319465909e-05,  \
+ 5.220102539170e-05, + 5.342696385924e-05, + 5.463024390338e-05, + 5.581025070569e-05, + 5.696639782400e-05,  \
+ 5.809849135403e-05, + 5.920614348724e-05, + 6.028912721376e-05, + 6.134756076790e-05, + 6.238130699785e-05,  \
+ 6.339056453726e-05, + 6.437556039600e-05, + 6.533659252455e-05, + 6.627410075453e-05, + 6.718833574269e-05 ]

* Data table for Id-Vg at Vd = 0.66V
.param vg_data_vd0.66=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.66=[ \
+ 5.214100000000e-10, + 7.550400000000e-10, + 1.093300000000e-09, + 1.583100000000e-09, + 2.292100000000e-09,  \
+ 3.318200000000e-09, + 4.803100000000e-09, + 6.951000000000e-09, + 1.005630000000e-08, + 1.454250000000e-08,  \
+ 2.101670000000e-08, + 3.034550000000e-08, + 4.375840000000e-08, + 6.298380000000e-08, + 9.042150000000e-08,  \
+ 1.293460000000e-07, + 1.841200000000e-07, + 2.603720000000e-07, + 3.650700000000e-07, + 5.063940000000e-07,  \
+ 6.933490000000e-07, + 9.351060000000e-07, + 1.240200000000e-06, + 1.615700000000e-06, + 2.066800000000e-06,  \
+ 2.596100000000e-06, + 3.204400000000e-06, + 3.890200000000e-06, + 4.650500000000e-06, + 5.481400000000e-06,  \
+ 6.378200000000e-06, + 7.335800000000e-06, + 8.349200000000e-06, + 9.413400000000e-06, + 1.052370000000e-05,  \
+ 1.167570000000e-05, + 1.286520000000e-05, + 1.408840000000e-05, + 1.534180000000e-05, + 1.662220000000e-05,  \
+ 1.792650000000e-05, + 1.925190000000e-05, + 2.059580000000e-05, + 2.195580000000e-05, + 2.332950000000e-05,  \
+ 2.471480000000e-05, + 2.610950000000e-05, + 2.751180000000e-05, + 2.891960000000e-05, + 3.033120000000e-05,  \
+ 3.174470000000e-05, + 3.315860000000e-05, + 3.457120000000e-05, + 3.598080000000e-05, + 3.738590000000e-05,  \
+ 3.878500000000e-05, + 4.017660000000e-05, + 4.155930000000e-05, + 4.293180000000e-05, + 4.429250000000e-05,  \
+ 4.564030000000e-05, + 4.697370000000e-05, + 4.829160000000e-05, + 4.959270000000e-05, + 5.087580000000e-05,  \
+ 5.213980000000e-05, + 5.338360000000e-05, + 5.460600000000e-05, + 5.580610000000e-05, + 5.698290000000e-05,  \
+ 5.813540000000e-05, + 5.926280000000e-05, + 6.036420000000e-05, + 6.143880000000e-05, + 6.248580000000e-05,  \
+ 6.350470000000e-05, + 6.449470000000e-05, + 6.545540000000e-05, + 6.638610000000e-05, + 6.728650000000e-05 ]

.param id_pred_data_vd0.66=[ \
+ 5.258934687724e-10, + 7.492223574879e-10, + 1.086110721360e-09, + 1.585480573496e-09, + 2.312790639003e-09,  \
+ 3.358607738591e-09, + 4.854167041657e-09, + 6.994934871329e-09, + 1.007228316752e-08, + 1.451393991658e-08,  \
+ 2.093558158833e-08, + 3.021090194011e-08, + 4.356854802268e-08, + 6.272949562458e-08, + 9.008984449110e-08,  \
+ 1.289386329972e-07, + 1.836809497036e-07, + 2.600065425895e-07, + 3.649268808203e-07, + 5.066072958471e-07,  \
+ 6.939699801478e-07, + 9.360784702039e-07, + 1.241413556272e-06, + 1.617162529328e-06, + 2.068678340947e-06,  \
+ 2.599156960059e-06, + 3.209585374861e-06, + 3.898932327502e-06, + 4.664457901526e-06, + 5.502142412297e-06,  \
+ 6.407131204469e-06, + 7.374056694971e-06, + 8.397409637837e-06, + 9.471763623878e-06, + 1.059202179022e-05,  \
+ 1.175330457045e-05, + 1.295131765801e-05, + 1.418204647052e-05, + 1.544197464682e-05, + 1.672791477176e-05,  \
+ 1.803701077733e-05, + 1.936663589731e-05, + 2.071443108434e-05, + 2.207819576142e-05, + 2.345590102777e-05,  \
+ 2.484546756023e-05, + 2.624507294968e-05, + 2.765275312413e-05, + 2.906671928940e-05, + 3.048505539482e-05,  \
+ 3.190589341102e-05, + 3.332747815875e-05, + 3.474792240013e-05, + 3.616535570472e-05, + 3.757805650821e-05,  \
+ 3.898417598975e-05, + 4.038201659569e-05, + 4.176986636594e-05, + 4.314595091273e-05, + 4.450893044122e-05,  \
+ 4.585711460095e-05, + 4.718921161839e-05, + 4.850382407312e-05, + 4.979983787052e-05, + 5.107589400723e-05,  \
+ 5.233147385297e-05, + 5.356517518521e-05, + 5.477647937369e-05, + 5.596471411991e-05, + 5.712923593819e-05,  \
+ 5.826979031553e-05, + 5.938597387285e-05, + 6.047755610780e-05, + 6.154446018627e-05, + 6.258665729547e-05,  \
+ 6.360427229083e-05, + 6.459739161073e-05, + 6.556642823853e-05, + 6.651154544670e-05, + 6.743317542714e-05 ]

* Data table for Id-Vg at Vd = 0.67V
.param vg_data_vd0.67=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.67=[ \
+ 5.263110000000e-10, + 7.620400000000e-10, + 1.103300000000e-09, + 1.597300000000e-09, + 2.312400000000e-09,  \
+ 3.347300000000e-09, + 4.844500000000e-09, + 7.010000000000e-09, + 1.014030000000e-08, + 1.466190000000e-08,  \
+ 2.118630000000e-08, + 3.058600000000e-08, + 4.409850000000e-08, + 6.346310000000e-08, + 9.109400000000e-08,  \
+ 1.302840000000e-07, + 1.854160000000e-07, + 2.621450000000e-07, + 3.674630000000e-07, + 5.095720000000e-07,  \
+ 6.974910000000e-07, + 9.403950000000e-07, + 1.246800000000e-06, + 1.623800000000e-06, + 2.076500000000e-06,  \
+ 2.607500000000e-06, + 3.217600000000e-06, + 3.905200000000e-06, + 4.667400000000e-06, + 5.500100000000e-06,  \
+ 6.398800000000e-06, + 7.358200000000e-06, + 8.373500000000e-06, + 9.439500000000e-06, + 1.055160000000e-05,  \
+ 1.170540000000e-05, + 1.289670000000e-05, + 1.412180000000e-05, + 1.537700000000e-05, + 1.665930000000e-05,  \
+ 1.796550000000e-05, + 1.929280000000e-05, + 2.063870000000e-05, + 2.200070000000e-05, + 2.337640000000e-05,  \
+ 2.476380000000e-05, + 2.616070000000e-05, + 2.756520000000e-05, + 2.897530000000e-05, + 3.038920000000e-05,  \
+ 3.180530000000e-05, + 3.322170000000e-05, + 3.463690000000e-05, + 3.604930000000e-05, + 3.745720000000e-05,  \
+ 3.885930000000e-05, + 4.025410000000e-05, + 4.164000000000e-05, + 4.301580000000e-05, + 4.438000000000e-05,  \
+ 4.573140000000e-05, + 4.706860000000e-05, + 4.839040000000e-05, + 4.969550000000e-05, + 5.098290000000e-05,  \
+ 5.225120000000e-05, + 5.349950000000e-05, + 5.472650000000e-05, + 5.593140000000e-05, + 5.711310000000e-05,  \
+ 5.827070000000e-05, + 5.940320000000e-05, + 6.050990000000e-05, + 6.158980000000e-05, + 6.264240000000e-05,  \
+ 6.366680000000e-05, + 6.466250000000e-05, + 6.562890000000e-05, + 6.656540000000e-05, + 6.747160000000e-05 ]

.param id_pred_data_vd0.67=[ \
+ 5.309481165838e-10, + 7.560067527557e-10, + 1.095523508576e-09, + 1.598919219248e-09, + 2.332318453924e-09,  \
+ 3.387153175716e-09, + 4.895694094564e-09, + 7.054749486812e-09, + 1.015752099320e-08, + 1.463442101723e-08,  \
+ 2.110550518353e-08, + 3.045064620011e-08, + 4.390834860146e-08, + 6.321295266787e-08, + 9.077732741503e-08,  \
+ 1.299116622988e-07, + 1.850438013662e-07, + 2.618862416170e-07, + 3.674690623257e-07, + 5.099725410673e-07,  \
+ 6.983253274484e-07, + 9.415895783604e-07, + 1.248237703066e-06, + 1.625446075195e-06, + 2.078550949136e-06,  \
+ 2.610741798890e-06, + 3.222996801924e-06, + 3.914257345059e-06, + 4.681795621764e-06, + 5.521566690732e-06,  \
+ 6.428665801650e-06, + 7.397761346510e-06, + 8.423287417827e-06, + 9.499792668066e-06, + 1.062212921170e-05,  \
+ 1.178547699965e-05, + 1.298540719290e-05, + 1.421797844159e-05, + 1.547959307572e-05, + 1.676711532127e-05,  \
+ 1.807760683732e-05, + 1.940857655427e-05, + 2.075762724417e-05, + 2.212258958025e-05, + 2.350140635826e-05,  \
+ 2.489212762157e-05, + 2.629288141179e-05, + 2.770183233224e-05, + 2.911711329944e-05, + 3.053697666473e-05,  \
+ 3.195953340764e-05, + 3.338309437822e-05, + 3.480580955511e-05, + 3.622581185482e-05, + 3.764148281334e-05,  \
+ 3.905087003659e-05, + 4.045233556099e-05, + 4.184431454632e-05, + 4.322504471929e-05, + 4.459294417757e-05,  \
+ 4.594651632942e-05, + 4.728450832772e-05, + 4.860538458161e-05, + 4.990797024220e-05, + 5.119119283336e-05,  \
+ 5.245390675555e-05, + 5.369530765165e-05, + 5.491447904205e-05, + 5.611084568955e-05, + 5.728375923354e-05,  \
+ 5.843274680956e-05, + 5.955744767562e-05, + 6.065767658583e-05, + 6.173317517096e-05, + 6.278395805566e-05,  \
+ 6.381001549016e-05, + 6.481160096882e-05, + 6.578886561329e-05, + 6.674202879367e-05, + 6.767149512598e-05 ]

* Data table for Id-Vg at Vd = 0.68V
.param vg_data_vd0.68=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.68=[ \
+ 5.312510000000e-10, + 7.690930000000e-10, + 1.113400000000e-09, + 1.611700000000e-09, + 2.332900000000e-09,  \
+ 3.376500000000e-09, + 4.886200000000e-09, + 7.069300000000e-09, + 1.022480000000e-08, + 1.478210000000e-08,  \
+ 2.135700000000e-08, + 3.082790000000e-08, + 4.444060000000e-08, + 6.394520000000e-08, + 9.177010000000e-08,  \
+ 1.312260000000e-07, + 1.867190000000e-07, + 2.639260000000e-07, + 3.698660000000e-07, + 5.127620000000e-07,  \
+ 7.016460000000e-07, + 9.456980000000e-07, + 1.253400000000e-06, + 1.631900000000e-06, + 2.086200000000e-06,  \
+ 2.618900000000e-06, + 3.230800000000e-06, + 3.920200000000e-06, + 4.684200000000e-06, + 5.518800000000e-06,  \
+ 6.419300000000e-06, + 7.380600000000e-06, + 8.397600000000e-06, + 9.465500000000e-06, + 1.057940000000e-05,  \
+ 1.173500000000e-05, + 1.292810000000e-05, + 1.415500000000e-05, + 1.541210000000e-05, + 1.669620000000e-05,  \
+ 1.800420000000e-05, + 1.933340000000e-05, + 2.068120000000e-05, + 2.204520000000e-05, + 2.342290000000e-05,  \
+ 2.481240000000e-05, + 2.621140000000e-05, + 2.761800000000e-05, + 2.903030000000e-05, + 3.044660000000e-05,  \
+ 3.186500000000e-05, + 3.328390000000e-05, + 3.470170000000e-05, + 3.611670000000e-05, + 3.752740000000e-05,  \
+ 3.893240000000e-05, + 4.033010000000e-05, + 4.171920000000e-05, + 4.309820000000e-05, + 4.446580000000e-05,  \
+ 4.582060000000e-05, + 4.716150000000e-05, + 4.848700000000e-05, + 4.979600000000e-05, + 5.108740000000e-05,  \
+ 5.235990000000e-05, + 5.361240000000e-05, + 5.484390000000e-05, + 5.605340000000e-05, + 5.723980000000e-05,  \
+ 5.840220000000e-05, + 5.953960000000e-05, + 6.065140000000e-05, + 6.173650000000e-05, + 6.279430000000e-05,  \
+ 6.382410000000e-05, + 6.482520000000e-05, + 6.579700000000e-05, + 6.673910000000e-05, + 6.765080000000e-05 ]

.param id_pred_data_vd0.68=[ \
+ 5.360546695421e-10, + 7.628251985636e-10, + 1.104942413122e-09, + 1.612309485921e-09, + 2.351720462812e-09,  \
+ 3.415466824919e-09, + 4.936890700691e-09, + 7.114141382658e-09, + 1.024229263180e-08, + 1.475447199084e-08,  \
+ 2.127490731141e-08, + 3.069014013590e-08, + 4.424820218674e-08, + 6.369687298502e-08, + 9.146642526048e-08,  \
+ 1.308878410100e-07, + 1.864114938144e-07, + 2.637720785970e-07, + 3.700192155520e-07, + 5.133446688887e-07,  \
+ 7.026842058622e-07, + 9.470937675360e-07, + 1.255037664123e-06, + 1.633679166844e-06, + 2.088344035656e-06,  \
+ 2.622201936902e-06, + 3.236224620196e-06, + 3.929351278202e-06, + 4.698823286162e-06, + 5.540602433030e-06,  \
+ 6.449764259742e-06, + 7.420929432556e-06, + 8.448554726783e-06, + 9.527135262033e-06, + 1.065150383511e-05,  \
+ 1.181680680020e-05, + 1.301861106185e-05, + 1.425292015483e-05, + 1.551615445351e-05, + 1.680514622421e-05,  \
+ 1.811705551518e-05, + 1.944926130818e-05, + 2.079941594275e-05, + 2.216543274699e-05, + 2.354521391680e-05,  \
+ 2.493688429240e-05, + 2.633860087371e-05, + 2.774854539894e-05, + 2.916499113780e-05, + 3.058610745938e-05,  \
+ 3.201009836630e-05, + 3.343530639540e-05, + 3.485988112516e-05, + 3.628215767094e-05, + 3.770039198571e-05,  \
+ 3.911273117410e-05, + 4.051761425217e-05, + 4.191327985609e-05, + 4.329818184488e-05, + 4.467065533390e-05,  \
+ 4.602939909091e-05, + 4.737273586215e-05, + 4.869951779256e-05, + 5.000843870221e-05, + 5.129840516020e-05,  \
+ 5.256817530608e-05, + 5.381699709687e-05, + 5.504397006007e-05, + 5.624836194329e-05, + 5.742946523242e-05,  \
+ 5.858690390596e-05, + 5.972021288471e-05, + 6.082901614718e-05, + 6.191316031618e-05, + 6.297265528701e-05,  \
+ 6.400753074558e-05, + 6.501761352411e-05, + 6.600326974876e-05, + 6.696477648802e-05, + 6.790226732846e-05 ]

* Data table for Id-Vg at Vd = 0.69V
.param vg_data_vd0.69=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.69=[ \
+ 5.362290000000e-10, + 7.762000000000e-10, + 1.123500000000e-09, + 1.626200000000e-09, + 2.353600000000e-09,  \
+ 3.405900000000e-09, + 4.928100000000e-09, + 7.129100000000e-09, + 1.030980000000e-08, + 1.490300000000e-08,  \
+ 2.152870000000e-08, + 3.107130000000e-08, + 4.478460000000e-08, + 6.442990000000e-08, + 9.244980000000e-08,  \
+ 1.321730000000e-07, + 1.880270000000e-07, + 2.657150000000e-07, + 3.722780000000e-07, + 5.159620000000e-07,  \
+ 7.058140000000e-07, + 9.510150000000e-07, + 1.260100000000e-06, + 1.640000000000e-06, + 2.095900000000e-06,  \
+ 2.630400000000e-06, + 3.243900000000e-06, + 3.935100000000e-06, + 4.701000000000e-06, + 5.537500000000e-06,  \
+ 6.439800000000e-06, + 7.402900000000e-06, + 8.421800000000e-06, + 9.491400000000e-06, + 1.060710000000e-05,  \
+ 1.176450000000e-05, + 1.295940000000e-05, + 1.418810000000e-05, + 1.544700000000e-05, + 1.673280000000e-05,  \
+ 1.804270000000e-05, + 1.937380000000e-05, + 2.072350000000e-05, + 2.208930000000e-05, + 2.346910000000e-05,  \
+ 2.486050000000e-05, + 2.626150000000e-05, + 2.767030000000e-05, + 2.908480000000e-05, + 3.050330000000e-05,  \
+ 3.192400000000e-05, + 3.334530000000e-05, + 3.476560000000e-05, + 3.618320000000e-05, + 3.759660000000e-05,  \
+ 3.900430000000e-05, + 4.040490000000e-05, + 4.179700000000e-05, + 4.317910000000e-05, + 4.454990000000e-05,  \
+ 4.590810000000e-05, + 4.725240000000e-05, + 4.858150000000e-05, + 4.989430000000e-05, + 5.118950000000e-05,  \
+ 5.246600000000e-05, + 5.372270000000e-05, + 5.495840000000e-05, + 5.617220000000e-05, + 5.736310000000e-05,  \
+ 5.853010000000e-05, + 5.967230000000e-05, + 6.078890000000e-05, + 6.187900000000e-05, + 6.294180000000e-05,  \
+ 6.397670000000e-05, + 6.498300000000e-05, + 6.596010000000e-05, + 6.690740000000e-05, + 6.782450000000e-05 ]

.param id_pred_data_vd0.69=[ \
+ 5.412171094621e-10, + 7.696854420480e-10, + 1.114367098598e-09, + 1.625636825153e-09, + 2.370978913202e-09,  \
+ 3.443535097070e-09, + 4.977737262379e-09, + 7.173084073386e-09, + 1.032648361488e-08, + 1.487387999433e-08,  \
+ 2.144364760426e-08, + 3.092901508239e-08, + 4.458767499216e-08, + 6.418077909132e-08, + 9.215628750781e-08,  \
+ 1.318657264449e-07, + 1.877825221186e-07, + 2.656627029296e-07, + 3.725732716475e-07, + 5.167204818690e-07,  \
+ 7.070387232488e-07, + 9.525821496936e-07, + 1.261803917032e-06, + 1.641852384182e-06, + 2.098037498399e-06,  \
+ 2.633514509398e-06, + 3.249246865380e-06, + 3.944162081098e-06, + 4.715500185739e-06, + 5.559211904256e-06,  \
+ 6.470341149907e-06, + 7.443510748999e-06, + 8.473148673147e-06, + 9.553748159306e-06, + 1.068005534762e-05,  \
+ 1.184723934784e-05, + 1.305083011175e-05, + 1.428680503523e-05, + 1.555160464704e-05, + 1.684203220066e-05,  \
+ 1.815517585783e-05, + 1.948852917849e-05, + 2.083969993691e-05, + 2.220660466264e-05, + 2.358724021178e-05,  \
+ 2.497970384866e-05, + 2.638221583766e-05, + 2.779295879009e-05, + 2.921024835814e-05, + 3.063234496949e-05,  \
+ 3.205757180694e-05, + 3.348412654304e-05, + 3.491031478916e-05, + 3.633451244241e-05, + 3.775489960390e-05,  \
+ 3.916983961972e-05, + 4.057770587679e-05, + 4.197676131298e-05, + 4.336545462138e-05, + 4.474215165828e-05,  \
+ 4.610557472915e-05, + 4.745408215967e-05, + 4.878639374510e-05, + 5.010132968891e-05, + 5.139761480677e-05,  \
+ 5.267426007777e-05, + 5.393023129727e-05, + 5.516468001588e-05, + 5.637681802909e-05, + 5.756605292845e-05,  \
+ 5.873179230548e-05, + 5.987361444568e-05, + 6.099107755290e-05, + 6.208403603523e-05, + 6.315228907624e-05,  \
+ 6.419581659429e-05, + 6.521471397718e-05, + 6.620898122492e-05, + 6.717905511323e-05, + 6.812487539719e-05 ]

* Data table for Id-Vg at Vd = 0.70V
.param vg_data_vd0.70=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.70=[ \
+ 5.412450000000e-10, + 7.833610000000e-10, + 1.133700000000e-09, + 1.640800000000e-09, + 2.374400000000e-09,  \
+ 3.435600000000e-09, + 4.970400000000e-09, + 7.189300000000e-09, + 1.039550000000e-08, + 1.502480000000e-08,  \
+ 2.170150000000e-08, + 3.131620000000e-08, + 4.513070000000e-08, + 6.491730000000e-08, + 9.313320000000e-08,  \
+ 1.331250000000e-07, + 1.893420000000e-07, + 2.675120000000e-07, + 3.747010000000e-07, + 5.191750000000e-07,  \
+ 7.099950000000e-07, + 9.563460000000e-07, + 1.266700000000e-06, + 1.648100000000e-06, + 2.105600000000e-06,  \
+ 2.641800000000e-06, + 3.257100000000e-06, + 3.950100000000e-06, + 4.717800000000e-06, + 5.556100000000e-06,  \
+ 6.460200000000e-06, + 7.425100000000e-06, + 8.445800000000e-06, + 9.517300000000e-06, + 1.063480000000e-05,  \
+ 1.179390000000e-05, + 1.299060000000e-05, + 1.422100000000e-05, + 1.548160000000e-05, + 1.676930000000e-05,  \
+ 1.808100000000e-05, + 1.941390000000e-05, + 2.076540000000e-05, + 2.213310000000e-05, + 2.351480000000e-05,  \
+ 2.490820000000e-05, + 2.631120000000e-05, + 2.772200000000e-05, + 2.913870000000e-05, + 3.055930000000e-05,  \
+ 3.198230000000e-05, + 3.340600000000e-05, + 3.482860000000e-05, + 3.624870000000e-05, + 3.766470000000e-05,  \
+ 3.907510000000e-05, + 4.047850000000e-05, + 4.187350000000e-05, + 4.325860000000e-05, + 4.463250000000e-05,  \
+ 4.599390000000e-05, + 4.734150000000e-05, + 4.867410000000e-05, + 4.999050000000e-05, + 5.128940000000e-05,  \
+ 5.256970000000e-05, + 5.383030000000e-05, + 5.507010000000e-05, + 5.628820000000e-05, + 5.748330000000e-05,  \
+ 5.865480000000e-05, + 5.980150000000e-05, + 6.092270000000e-05, + 6.201750000000e-05, + 6.308510000000e-05,  \
+ 6.412490000000e-05, + 6.513620000000e-05, + 6.611830000000e-05, + 6.707070000000e-05, + 6.799290000000e-05 ]

.param id_pred_data_vd0.70=[ \
+ 5.464385166576e-10, + 7.765894149969e-10, + 1.123796811164e-09, + 1.638905211543e-09, + 2.390084574699e-09,  \
+ 3.471336285088e-09, + 5.018193105499e-09, + 7.231520360307e-09, + 1.041009198843e-08, + 1.499253396986e-08,  \
+ 2.161166214876e-08, + 3.116706643880e-08, + 4.492639789078e-08, + 6.466415385376e-08, + 9.284618727179e-08,  \
+ 1.328444156456e-07, + 1.891545764465e-07, + 2.675548017805e-07, + 3.751284282316e-07, + 5.200925500048e-07,  \
+ 7.113833930816e-07, + 9.580491337147e-07, + 1.268522748887e-06, + 1.649945102145e-06, + 2.107608634105e-06,  \
+ 2.644653204698e-06, + 3.262031395934e-06, + 3.958669185522e-06, + 4.731788249046e-06, + 5.577334104601e-06,  \
+ 6.490362557088e-06, + 7.465454473277e-06, + 8.497000999341e-06, + 9.579518700775e-06, + 1.070771068044e-05,  \
+ 1.187669258798e-05, + 1.308199134655e-05, + 1.431959353795e-05, + 1.558583844599e-05, + 1.687759249762e-05,  \
+ 1.819192966650e-05, + 1.952632628672e-05, + 2.087842549372e-05, + 2.224610980193e-05, + 2.362744126003e-05,  \
+ 2.502051502233e-05, + 2.642362742336e-05, + 2.783501877275e-05, + 2.925294975284e-05, + 3.067577781621e-05,  \
+ 3.210192408005e-05, + 3.352952444402e-05, + 3.495707896946e-05, + 3.638280250016e-05, + 3.780511360674e-05,  \
+ 3.922227297153e-05, + 4.063268133905e-05, + 4.203471653454e-05, + 4.342682004790e-05, + 4.480742572923e-05,  \
+ 4.617504382622e-05, + 4.752829918289e-05, + 4.886586757493e-05, + 5.018638912588e-05, + 5.148874843144e-05,  \
+ 5.277188611217e-05, + 5.403477844084e-05, + 5.527641187655e-05, + 5.649623126374e-05, + 5.769332492491e-05,  \
+ 5.886719882255e-05, + 6.001737419865e-05, + 6.114329589764e-05, + 6.224509124877e-05, + 6.332215925795e-05,  \
+ 6.437450501835e-05, + 6.540229151142e-05, + 6.640543215326e-05, + 6.738410520484e-05, + 6.833874358563e-05 ]

* Data table for Id-Vg at Vd = 0.71V
.param vg_data_vd0.71=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.71=[ \
+ 5.463010000000e-10, + 7.905770000000e-10, + 1.144000000000e-09, + 1.655500000000e-09, + 2.395300000000e-09,  \
+ 3.465400000000e-09, + 5.012900000000e-09, + 7.249800000000e-09, + 1.048170000000e-08, + 1.514730000000e-08,  \
+ 2.187540000000e-08, + 3.156250000000e-08, + 4.547880000000e-08, + 6.540760000000e-08, + 9.382020000000e-08,  \
+ 1.340820000000e-07, + 1.906640000000e-07, + 2.693170000000e-07, + 3.771330000000e-07, + 5.223990000000e-07,  \
+ 7.141890000000e-07, + 9.616920000000e-07, + 1.273400000000e-06, + 1.656300000000e-06, + 2.115300000000e-06,  \
+ 2.653200000000e-06, + 3.270300000000e-06, + 3.965100000000e-06, + 4.734600000000e-06, + 5.574700000000e-06,  \
+ 6.480600000000e-06, + 7.447400000000e-06, + 8.469800000000e-06, + 9.543000000000e-06, + 1.066230000000e-05,  \
+ 1.182320000000e-05, + 1.302160000000e-05, + 1.425380000000e-05, + 1.551620000000e-05, + 1.680560000000e-05,  \
+ 1.811900000000e-05, + 1.945370000000e-05, + 2.080700000000e-05, + 2.217660000000e-05, + 2.356010000000e-05,  \
+ 2.495540000000e-05, + 2.636050000000e-05, + 2.777330000000e-05, + 2.919200000000e-05, + 3.061480000000e-05,  \
+ 3.204000000000e-05, + 3.346590000000e-05, + 3.489090000000e-05, + 3.631340000000e-05, + 3.773190000000e-05,  \
+ 3.914490000000e-05, + 4.055100000000e-05, + 4.194870000000e-05, + 4.333670000000e-05, + 4.471360000000e-05,  \
+ 4.607810000000e-05, + 4.742900000000e-05, + 4.876490000000e-05, + 5.008470000000e-05, + 5.138710000000e-05,  \
+ 5.267110000000e-05, + 5.393550000000e-05, + 5.517920000000e-05, + 5.640130000000e-05, + 5.760060000000e-05,  \
+ 5.877620000000e-05, + 5.992730000000e-05, + 6.105290000000e-05, + 6.215230000000e-05, + 6.322450000000e-05,  \
+ 6.426900000000e-05, + 6.528510000000e-05, + 6.627200000000e-05, + 6.722930000000e-05, + 6.815640000000e-05 ]

.param id_pred_data_vd0.71=[ \
+ 5.517197532168e-10, + 7.835373894149e-10, + 1.133230705941e-09, + 1.652121233153e-09, + 2.409027077821e-09,  \
+ 3.498861560480e-09, + 5.058234582300e-09, + 7.289389429843e-09, + 1.049295711653e-08, + 1.511037650559e-08,  \
+ 2.177862214126e-08, + 3.140407383029e-08, + 4.526389297155e-08, + 6.514669451008e-08, + 9.353537620882e-08,  \
+ 1.338227180270e-07, + 1.905268402425e-07, + 2.694462267527e-07, + 3.776812565093e-07, + 5.234571796109e-07,  \
+ 7.157104494127e-07, + 9.634785374146e-07, + 1.275187438523e-06, + 1.657947893818e-06, + 2.117037788594e-06,  \
+ 2.655590662926e-06, + 3.274548007539e-06, + 3.972827721554e-06, + 4.747647790282e-06, + 5.594944886980e-06,  \
+ 6.509769727927e-06, + 7.486684526157e-06, + 8.520075853085e-06, + 9.604415517970e-06, + 1.073438196727e-05,  \
+ 1.190509598018e-05, + 1.311202639044e-05, + 1.435114183550e-05, + 1.561883649629e-05, + 1.691180934358e-05,  \
+ 1.822722944780e-05, + 1.956255387995e-05, + 2.091546572046e-05, + 2.228385597846e-05, + 2.366574997723e-05,  \
+ 2.505931122869e-05, + 2.646288405231e-05, + 2.787464487483e-05, + 2.929305683210e-05, + 3.071645907767e-05,  \
+ 3.214314685465e-05, + 3.357158846484e-05, + 3.500013339362e-05, + 3.642712596047e-05, + 3.785099055676e-05,  \
+ 3.927001984266e-05, + 4.068260979693e-05, + 4.208729071252e-05, + 4.348233458586e-05, + 4.486638019443e-05,  \
+ 4.623795524822e-05, + 4.759555129567e-05, + 4.893790268397e-05, + 5.026372826251e-05, + 5.157183470146e-05,  \
+ 5.286102867103e-05, + 5.413048878836e-05, + 5.537907338294e-05, + 5.660623486619e-05, + 5.781095038401e-05,  \
+ 5.899278599827e-05, + 6.015120961820e-05, + 6.128566332336e-05, + 6.239603346330e-05, + 6.348188609991e-05,  \
+ 6.454316440795e-05, + 6.557977023476e-05, + 6.659185855824e-05, + 6.757959985407e-05, + 6.854281848064e-05 ]

* Data table for Id-Vg at Vd = 0.72V
.param vg_data_vd0.72=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.72=[ \
+ 5.513960000000e-10, + 7.978480000000e-10, + 1.154400000000e-09, + 1.670200000000e-09, + 2.416400000000e-09,  \
+ 3.495500000000e-09, + 5.055800000000e-09, + 7.310800000000e-09, + 1.056840000000e-08, + 1.527060000000e-08,  \
+ 2.205030000000e-08, + 3.181030000000e-08, + 4.582900000000e-08, + 6.590060000000e-08, + 9.451100000000e-08,  \
+ 1.350440000000e-07, + 1.919920000000e-07, + 2.711300000000e-07, + 3.795750000000e-07, + 5.256360000000e-07,  \
+ 7.183980000000e-07, + 9.670520000000e-07, + 1.280100000000e-06, + 1.664400000000e-06, + 2.125100000000e-06,  \
+ 2.664600000000e-06, + 3.283500000000e-06, + 3.980100000000e-06, + 4.751400000000e-06, + 5.593300000000e-06,  \
+ 6.501000000000e-06, + 7.469500000000e-06, + 8.493800000000e-06, + 9.568700000000e-06, + 1.068970000000e-05,  \
+ 1.185230000000e-05, + 1.305250000000e-05, + 1.428640000000e-05, + 1.555050000000e-05, + 1.684170000000e-05,  \
+ 1.815680000000e-05, + 1.949330000000e-05, + 2.084840000000e-05, + 2.221980000000e-05, + 2.360510000000e-05,  \
+ 2.500230000000e-05, + 2.640930000000e-05, + 2.782400000000e-05, + 2.924480000000e-05, + 3.066960000000e-05,  \
+ 3.209700000000e-05, + 3.352510000000e-05, + 3.495230000000e-05, + 3.637720000000e-05, + 3.779810000000e-05,  \
+ 3.921360000000e-05, + 4.062230000000e-05, + 4.202270000000e-05, + 4.341350000000e-05, + 4.479330000000e-05,  \
+ 4.616080000000e-05, + 4.751470000000e-05, + 4.885390000000e-05, + 5.017700000000e-05, + 5.148280000000e-05,  \
+ 5.277040000000e-05, + 5.403840000000e-05, + 5.528590000000e-05, + 5.651180000000e-05, + 5.771500000000e-05,  \
+ 5.889480000000e-05, + 6.005000000000e-05, + 6.117980000000e-05, + 6.228350000000e-05, + 6.336020000000e-05,  \
+ 6.440920000000e-05, + 6.542980000000e-05, + 6.642140000000e-05, + 6.738340000000e-05, + 6.831520000000e-05 ]

.param id_pred_data_vd0.72=[ \
+ 5.570626759877e-10, + 7.905324395097e-10, + 1.142678272004e-09, + 1.665272080231e-09, + 2.427813949879e-09,  \
+ 3.526093976802e-09, + 5.097817528110e-09, + 7.346628265736e-09, + 1.057502885260e-08, + 1.522722811842e-08,  \
+ 2.194444562065e-08, + 3.163968415265e-08, + 4.560000888887e-08, + 6.562757505435e-08, + 9.422275184079e-08,  \
+ 1.347994714251e-07, + 1.918969815051e-07, + 2.713344633776e-07, + 3.802282571996e-07, + 5.268098584565e-07,  \
+ 7.200149775599e-07, + 9.688703266875e-07, + 1.281778313569e-06, + 1.665840063652e-06, + 2.126314157067e-06,  \
+ 2.666314012458e-06, + 3.286773753644e-06, + 3.986607334809e-06, + 4.763038086821e-06, + 5.611984088318e-06,  \
+ 6.528505909955e-06, + 7.507144182455e-06, + 8.542267969460e-06, + 9.628320331103e-06, + 1.076000167814e-05,  \
+ 1.193236079416e-05, + 1.314084001933e-05, + 1.438141538529e-05, + 1.565041064168e-05, + 1.694455946563e-05,  \
+ 1.826102903578e-05, + 1.959720393643e-05, + 2.095083415043e-05, + 2.231979276985e-05, + 2.370212838287e-05,  \
+ 2.509606245439e-05, + 2.649984788150e-05, + 2.791190257994e-05, + 2.933056064649e-05, + 3.075426095165e-05,  \
+ 3.218138474040e-05, + 3.361030801898e-05, + 3.503963205731e-05, + 3.646750235930e-05, + 3.789258567849e-05,  \
+ 3.931313491194e-05, + 4.072758631082e-05, + 4.213446256472e-05, + 4.353219468612e-05, + 4.491932108067e-05,  \
+ 4.629432514776e-05, + 4.765585006680e-05, + 4.900261759758e-05, + 5.033326568082e-05, + 5.164667847566e-05,  \
+ 5.294178205077e-05, + 5.421736626886e-05, + 5.547266628128e-05, + 5.670677055605e-05, + 5.791881470941e-05,  \
+ 5.910849489737e-05, + 6.027482100762e-05, + 6.141769874375e-05, + 6.253648374695e-05, + 6.363109219819e-05,  \
+ 6.470115738921e-05, + 6.574682076462e-05, + 6.676791992504e-05, + 6.776460155379e-05, + 6.873688660562e-05 ]

* Data table for Id-Vg at Vd = 0.73V
.param vg_data_vd0.73=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.73=[ \
+ 5.565310000000e-10, + 8.051750000000e-10, + 1.164900000000e-09, + 1.685200000000e-09, + 2.437600000000e-09,  \
+ 3.525800000000e-09, + 5.098900000000e-09, + 7.372200000000e-09, + 1.065570000000e-08, + 1.539460000000e-08,  \
+ 2.222640000000e-08, + 3.205970000000e-08, + 4.618120000000e-08, + 6.639630000000e-08, + 9.520560000000e-08,  \
+ 1.360110000000e-07, + 1.933260000000e-07, + 2.729520000000e-07, + 3.820280000000e-07, + 5.288840000000e-07,  \
+ 7.226190000000e-07, + 9.724270000000e-07, + 1.286800000000e-06, + 1.672600000000e-06, + 2.134900000000e-06,  \
+ 2.676100000000e-06, + 3.296700000000e-06, + 3.995000000000e-06, + 4.768100000000e-06, + 5.611800000000e-06,  \
+ 6.521400000000e-06, + 7.491700000000e-06, + 8.517600000000e-06, + 9.594400000000e-06, + 1.071710000000e-05,  \
+ 1.188140000000e-05, + 1.308330000000e-05, + 1.431890000000e-05, + 1.558470000000e-05, + 1.687750000000e-05,  \
+ 1.819440000000e-05, + 1.953260000000e-05, + 2.088950000000e-05, + 2.226270000000e-05, + 2.364980000000e-05,  \
+ 2.504880000000e-05, + 2.645770000000e-05, + 2.787440000000e-05, + 2.929700000000e-05, + 3.072400000000e-05,  \
+ 3.215340000000e-05, + 3.358360000000e-05, + 3.501310000000e-05, + 3.644020000000e-05, + 3.786350000000e-05,  \
+ 3.928140000000e-05, + 4.069260000000e-05, + 4.209560000000e-05, + 4.348910000000e-05, + 4.487170000000e-05,  \
+ 4.624210000000e-05, + 4.759900000000e-05, + 4.894120000000e-05, + 5.026750000000e-05, + 5.157670000000e-05,  \
+ 5.286760000000e-05, + 5.413910000000e-05, + 5.539020000000e-05, + 5.661980000000e-05, + 5.782680000000e-05,  \
+ 5.901050000000e-05, + 6.016970000000e-05, + 6.130360000000e-05, + 6.241150000000e-05, + 6.349240000000e-05,  \
+ 6.454570000000e-05, + 6.557070000000e-05, + 6.656670000000e-05, + 6.753320000000e-05, + 6.846960000000e-05 ]

.param id_pred_data_vd0.73=[ \
+ 5.624710763819e-10, + 7.975775839775e-10, + 1.152134071480e-09, + 1.678370409319e-09, + 2.446434017589e-09,  \
+ 3.553015135438e-09, + 5.136934695393e-09, + 7.403199102640e-09, + 1.065625546914e-08, + 1.534295959615e-08,  \
+ 2.210895338806e-08, + 3.187371014235e-08, + 4.593431398803e-08, + 6.610643502825e-08, + 9.490809432577e-08,  \
+ 1.357734808494e-07, + 1.932636510560e-07, + 2.732176199061e-07, + 3.827660492561e-07, + 5.301454820028e-07,  \
+ 7.242878666602e-07, + 9.742065662977e-07, + 1.288288566457e-06, + 1.673609879163e-06, + 2.135406680281e-06,  \
+ 2.676786250504e-06, + 3.298672781966e-06, + 3.999968298558e-06, + 4.777902713613e-06, + 5.628408453049e-06,  \
+ 6.546513668582e-06, + 7.526774788857e-06, + 8.563535120629e-06, + 9.651214986661e-06, + 1.078449696251e-05,  \
+ 1.195840621222e-05, + 1.316835563557e-05, + 1.441029193302e-05, + 1.568051966387e-05, + 1.697578158200e-05,  \
+ 1.829317763622e-05, + 1.963015036381e-05, + 2.098439459587e-05, + 2.235381762148e-05, + 2.373647279455e-05,  \
+ 2.513065381208e-05, + 2.653457868291e-05, + 2.794672567688e-05, + 2.936549870356e-05, + 3.078922200075e-05,  \
+ 3.221652521461e-05, + 3.364578835317e-05, + 3.507544985041e-05, + 3.650401718915e-05, + 3.792994473770e-05,  \
+ 3.935163374990e-05, + 4.076766606886e-05, + 4.217636858812e-05, + 4.357640282251e-05, + 4.496618596022e-05,  \
+ 4.634421486116e-05, + 4.770939005539e-05, + 4.906009686238e-05, + 5.039519332058e-05, + 5.171352684556e-05,  \
+ 5.301389173837e-05, + 5.429541160993e-05, + 5.555697105592e-05, + 5.679771493305e-05, + 5.801690494991e-05,  \
+ 5.921390373260e-05, + 6.038818544766e-05, + 6.153902242659e-05, + 6.266623408010e-05, + 6.376943798386e-05,  \
+ 6.484832607384e-05, + 6.590290366148e-05, + 6.693300078041e-05, + 6.793875552830e-05, + 6.892017321661e-05 ]

* Data table for Id-Vg at Vd = 0.74V
.param vg_data_vd0.74=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.74=[ \
+ 5.617060000000e-10, + 8.125580000000e-10, + 1.175400000000e-09, + 1.700200000000e-09, + 2.459000000000e-09,  \
+ 3.556300000000e-09, + 5.142300000000e-09, + 7.434000000000e-09, + 1.074360000000e-08, + 1.551950000000e-08,  \
+ 2.240360000000e-08, + 3.231050000000e-08, + 4.653550000000e-08, + 6.689500000000e-08, + 9.590400000000e-08,  \
+ 1.369820000000e-07, + 1.946670000000e-07, + 2.747820000000e-07, + 3.844910000000e-07, + 5.321440000000e-07,  \
+ 7.268550000000e-07, + 9.778170000000e-07, + 1.293500000000e-06, + 1.680800000000e-06, + 2.144600000000e-06,  \
+ 2.687500000000e-06, + 3.309900000000e-06, + 4.010000000000e-06, + 4.784900000000e-06, + 5.630400000000e-06,  \
+ 6.541700000000e-06, + 7.513800000000e-06, + 8.541500000000e-06, + 9.619900000000e-06, + 1.074440000000e-05,  \
+ 1.191040000000e-05, + 1.311390000000e-05, + 1.435120000000e-05, + 1.561870000000e-05, + 1.691330000000e-05,  \
+ 1.823190000000e-05, + 1.957180000000e-05, + 2.093040000000e-05, + 2.230530000000e-05, + 2.369420000000e-05,  \
+ 2.509500000000e-05, + 2.650570000000e-05, + 2.792420000000e-05, + 2.934880000000e-05, + 3.077770000000e-05,  \
+ 3.220920000000e-05, + 3.364150000000e-05, + 3.507310000000e-05, + 3.650250000000e-05, + 3.792800000000e-05,  \
+ 3.934830000000e-05, + 4.076200000000e-05, + 4.216750000000e-05, + 4.356360000000e-05, + 4.494880000000e-05,  \
+ 4.632200000000e-05, + 4.768180000000e-05, + 4.902700000000e-05, + 5.035630000000e-05, + 5.166870000000e-05,  \
+ 5.296280000000e-05, + 5.423770000000e-05, + 5.549230000000e-05, + 5.672540000000e-05, + 5.793610000000e-05,  \
+ 5.912350000000e-05, + 6.028660000000e-05, + 6.142440000000e-05, + 6.253630000000e-05, + 6.362130000000e-05,  \
+ 6.467880000000e-05, + 6.570790000000e-05, + 6.670820000000e-05, + 6.767900000000e-05, + 6.861970000000e-05 ]

.param id_pred_data_vd0.74=[ \
+ 5.679467607322e-10, + 8.046725930022e-10, + 1.161600702293e-09, + 1.691402609083e-09, + 2.464884731879e-09,  \
+ 3.579620324601e-09, + 5.175548531966e-09, + 7.459089541584e-09, + 1.073650111039e-08, + 1.545749512388e-08,  \
+ 2.227195778914e-08, + 3.210601505543e-08, + 4.626635757177e-08, + 6.658239641411e-08, + 9.559005178517e-08,  \
+ 1.367433355881e-07, + 1.946248613649e-07, + 2.750924062411e-07, + 3.852896372791e-07, + 5.334570437299e-07,  \
+ 7.285244828381e-07, + 9.794854759093e-07, + 1.294704979955e-06, + 1.681238159108e-06, + 2.144303321074e-06,  \
+ 2.686984944376e-06, + 3.310214833618e-06, + 4.012888721263e-06, + 4.792225327037e-06, + 5.644160919474e-06,  \
+ 6.563752122020e-06, + 7.545515454694e-06, + 8.583784710936e-06, + 9.672993965069e-06, + 1.080777112293e-05,  \
+ 1.198312838824e-05, + 1.319447168498e-05, + 1.443770161131e-05, + 1.570907075802e-05, + 1.700536206044e-05,  \
+ 1.832360208937e-05, + 1.966129930224e-05, + 2.101606984070e-05, + 2.238589462650e-05, + 2.376878823270e-05,  \
+ 2.516306674806e-05, + 2.656700453372e-05, + 2.797911285597e-05, + 2.939768222859e-05, + 3.082140698098e-05,  \
+ 3.224863416108e-05, + 3.367794233782e-05, + 3.510779701173e-05, + 3.653673906229e-05, + 3.796322322160e-05,  \
+ 3.938581998227e-05, + 4.080296523171e-05, + 4.221308947308e-05, + 4.361496779893e-05, + 4.500696610194e-05,  \
+ 4.638774640625e-05, + 4.775602996233e-05, + 4.911030919175e-05, + 5.044946417911e-05, + 5.177237500902e-05,  \
+ 5.307771178195e-05, + 5.436461302452e-05, + 5.563213111600e-05, + 5.687916229363e-05, + 5.810519505758e-05,  \
+ 5.930933562922e-05, + 6.049105097190e-05, + 6.164978112793e-05, + 6.278519227635e-05, + 6.389676753315e-05,  \
+ 6.498431306682e-05, + 6.604759197216e-05, + 6.708679269650e-05, + 6.810154911363e-05, + 6.909197429195e-05 ]

* Data table for Id-Vg at Vd = 0.75V
.param vg_data_vd0.75=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.75=[ \
+ 5.669220000000e-10, + 8.199970000000e-10, + 1.186000000000e-09, + 1.715300000000e-09, + 2.480600000000e-09,  \
+ 3.587000000000e-09, + 5.186000000000e-09, + 7.496300000000e-09, + 1.083210000000e-08, + 1.564520000000e-08,  \
+ 2.258180000000e-08, + 3.256290000000e-08, + 4.689190000000e-08, + 6.739640000000e-08, + 9.660610000000e-08,  \
+ 1.379590000000e-07, + 1.960140000000e-07, + 2.766200000000e-07, + 3.869640000000e-07, + 5.354170000000e-07,  \
+ 7.311050000000e-07, + 9.832220000000e-07, + 1.300200000000e-06, + 1.689000000000e-06, + 2.154400000000e-06,  \
+ 2.699000000000e-06, + 3.323100000000e-06, + 4.025000000000e-06, + 4.801700000000e-06, + 5.648900000000e-06,  \
+ 6.562000000000e-06, + 7.535800000000e-06, + 8.565300000000e-06, + 9.645400000000e-06, + 1.077160000000e-05,  \
+ 1.193930000000e-05, + 1.314450000000e-05, + 1.438340000000e-05, + 1.565260000000e-05, + 1.694880000000e-05,  \
+ 1.826910000000e-05, + 1.961070000000e-05, + 2.097100000000e-05, + 2.234760000000e-05, + 2.373820000000e-05,  \
+ 2.514080000000e-05, + 2.655330000000e-05, + 2.797370000000e-05, + 2.940020000000e-05, + 3.083100000000e-05,  \
+ 3.226440000000e-05, + 3.369880000000e-05, + 3.513250000000e-05, + 3.656400000000e-05, + 3.799180000000e-05,  \
+ 3.941440000000e-05, + 4.083030000000e-05, + 4.223830000000e-05, + 4.363690000000e-05, + 4.502480000000e-05,  \
+ 4.640060000000e-05, + 4.776320000000e-05, + 4.911130000000e-05, + 5.044360000000e-05, + 5.175900000000e-05,  \
+ 5.305630000000e-05, + 5.433440000000e-05, + 5.559230000000e-05, + 5.682880000000e-05, + 5.804310000000e-05,  \
+ 5.923400000000e-05, + 6.040080000000e-05, + 6.154240000000e-05, + 6.265810000000e-05, + 6.374700000000e-05,  \
+ 6.480850000000e-05, + 6.584170000000e-05, + 6.684610000000e-05, + 6.782100000000e-05, + 6.876590000000e-05 ]

.param id_pred_data_vd0.75=[ \
+ 5.734935026869e-10, + 8.118217764697e-10, + 1.171085395324e-09, + 1.704374308353e-09, + 2.483153682675e-09,  \
+ 3.605889919989e-09, + 5.213639520107e-09, + 7.514216582294e-09, + 1.081578759887e-08, + 1.557075401948e-08,  \
+ 2.243330587959e-08, + 3.233607781539e-08, + 4.659584718070e-08, + 6.705541721885e-08, + 9.626804953200e-08,  \
+ 1.377082341492e-07, + 1.959793181072e-07, + 2.769566549432e-07, + 3.877967600374e-07, + 5.367424478209e-07,  \
+ 7.327155628900e-07, + 9.846901320998e-07, + 1.301012588328e-06, + 1.688710312919e-06, + 2.152979448056e-06,  \
+ 2.696897297483e-06, + 3.321368012621e-06, + 4.025315206491e-06, + 4.805951220987e-06, + 5.659220505549e-06,  \
+ 6.580154831681e-06, + 7.563289045720e-06, + 8.602978596173e-06, + 9.693597348814e-06, + 1.082975859390e-05,  \
+ 1.200645419885e-05, + 1.321910849583e-05, + 1.446351416234e-05, + 1.573600138727e-05, + 1.703321549940e-05,  \
+ 1.835228476921e-05, + 1.969059258045e-05, + 2.104583472828e-05, + 2.241593347208e-05, + 2.379900342930e-05,  \
+ 2.519325062167e-05, + 2.659707206476e-05, + 2.800893707899e-05, + 2.942730407085e-05, + 3.085072967224e-05,  \
+ 3.227768047509e-05, + 3.370683043613e-05, + 3.513660522003e-05, + 3.656563785626e-05, + 3.799241676461e-05,  \
+ 3.941554496123e-05, + 4.083344811079e-05, + 4.224486838211e-05, + 4.364813321445e-05, + 4.504209118750e-05,  \
+ 4.642505882657e-05, + 4.779599112226e-05, + 4.915355930279e-05, + 5.049630090070e-05, + 5.182326094655e-05,  \
+ 5.313327710610e-05, + 5.442520341603e-05, + 5.569817221840e-05, + 5.695124491467e-05, + 5.818360841658e-05,  \
+ 5.939458606008e-05, + 6.058348481019e-05, + 6.174975897011e-05, + 6.289294469752e-05, + 6.401277460100e-05,  \
+ 6.510875755339e-05, + 6.618088264077e-05, + 6.722878970322e-05, + 6.825258788012e-05, + 6.925234265509e-05 ]

* Data table for Id-Vg at Vd = 0.76V
.param vg_data_vd0.76=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.76=[ \
+ 5.721780000000e-10, + 8.274940000000e-10, + 1.196700000000e-09, + 1.730500000000e-09, + 2.502300000000e-09,  \
+ 3.617900000000e-09, + 5.230100000000e-09, + 7.558900000000e-09, + 1.092120000000e-08, + 1.577170000000e-08,  \
+ 2.276120000000e-08, + 3.281690000000e-08, + 4.725040000000e-08, + 6.790070000000e-08, + 9.731220000000e-08,  \
+ 1.389410000000e-07, + 1.973680000000e-07, + 2.784660000000e-07, + 3.894470000000e-07, + 5.387020000000e-07,  \
+ 7.353680000000e-07, + 9.886430000000e-07, + 1.307000000000e-06, + 1.697200000000e-06, + 2.164200000000e-06,  \
+ 2.710500000000e-06, + 3.336300000000e-06, + 4.040000000000e-06, + 4.818400000000e-06, + 5.667400000000e-06,  \
+ 6.582300000000e-06, + 7.557800000000e-06, + 8.589000000000e-06, + 9.670900000000e-06, + 1.079870000000e-05,  \
+ 1.196810000000e-05, + 1.317500000000e-05, + 1.441550000000e-05, + 1.568640000000e-05, + 1.698420000000e-05,  \
+ 1.830610000000e-05, + 1.964930000000e-05, + 2.101130000000e-05, + 2.238960000000e-05, + 2.378200000000e-05,  \
+ 2.518630000000e-05, + 2.660060000000e-05, + 2.802280000000e-05, + 2.945110000000e-05, + 3.088380000000e-05,  \
+ 3.231910000000e-05, + 3.375550000000e-05, + 3.519120000000e-05, + 3.662480000000e-05, + 3.805470000000e-05,  \
+ 3.947960000000e-05, + 4.089780000000e-05, + 4.230820000000e-05, + 4.370920000000e-05, + 4.509960000000e-05,  \
+ 4.647810000000e-05, + 4.784330000000e-05, + 4.919410000000e-05, + 5.052930000000e-05, + 5.184760000000e-05,  \
+ 5.314800000000e-05, + 5.442920000000e-05, + 5.569030000000e-05, + 5.693010000000e-05, + 5.814780000000e-05,  \
+ 5.934220000000e-05, + 6.051240000000e-05, + 6.165770000000e-05, + 6.277710000000e-05, + 6.386980000000e-05,  \
+ 6.493500000000e-05, + 6.597220000000e-05, + 6.698050000000e-05, + 6.795940000000e-05, + 6.890830000000e-05 ]

.param id_pred_data_vd0.76=[ \
+ 5.791107748898e-10, + 8.190295019972e-10, + 1.180581779003e-09, + 1.717290816217e-09, + 2.501256464171e-09,  \
+ 3.631831315687e-09, + 5.251187324973e-09, + 7.568549627024e-09, + 1.089397212439e-08, + 1.568259285989e-08,  \
+ 2.259284229922e-08, + 3.256398912299e-08, + 4.692238093185e-08, + 6.752481283456e-08, + 9.694138782379e-08,  \
+ 1.386666616554e-07, + 1.973241023734e-07, + 2.788071037685e-07, + 3.902827870661e-07, + 5.399958467933e-07,  \
+ 7.368538535957e-07, + 9.898182497636e-07, + 1.307203197030e-06, + 1.696012959655e-06, + 2.161421634810e-06,  \
+ 2.706483619477e-06, + 3.332112701173e-06, + 4.037220041937e-06, + 4.819043715543e-06, + 5.673495525116e-06,  \
+ 6.595664381166e-06, + 7.580060300825e-06, + 8.621027409390e-06, + 9.712933679111e-06, + 1.085037863959e-05,  \
+ 1.202833991556e-05, + 1.324218152149e-05, + 1.448770985007e-05, + 1.576118265803e-05, + 1.705926828436e-05,  \
+ 1.837905809225e-05, + 1.971790748939e-05, + 2.107354237523e-05, + 2.244383933430e-05, + 2.382697217399e-05,  \
+ 2.522112714360e-05, + 2.662472412339e-05, + 2.803626455716e-05, + 2.945424988866e-05, + 3.087723962381e-05,  \
+ 3.230375179555e-05, + 3.373254221515e-05, + 3.516200173181e-05, + 3.659088062705e-05, + 3.801766652032e-05,  \
+ 3.944091062294e-05, + 4.085937704076e-05, + 4.227156998240e-05, + 4.367601577542e-05, + 4.507138175541e-05,  \
+ 4.645639884984e-05, + 4.782962379977e-05, + 4.918978753267e-05, + 5.053588363808e-05, + 5.186645226786e-05,  \
+ 5.318055336829e-05, + 5.447716946946e-05, + 5.575522780418e-05, + 5.701383255655e-05, + 5.825220956467e-05,  \
+ 5.946960678557e-05, + 6.066532747354e-05, + 6.183890160173e-05, + 6.298974301899e-05, + 6.411747570382e-05,  \
+ 6.522171257529e-05, + 6.630221585510e-05, + 6.735891365679e-05, + 6.839167326689e-05, + 6.940035091247e-05 ]

* Data table for Id-Vg at Vd = 0.77V
.param vg_data_vd0.77=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.77=[ \
+ 5.774750000000e-10, + 8.350490000000e-10, + 1.207500000000e-09, + 1.745900000000e-09, + 2.524200000000e-09,  \
+ 3.649100000000e-09, + 5.274400000000e-09, + 7.622000000000e-09, + 1.101090000000e-08, + 1.589900000000e-08,  \
+ 2.294180000000e-08, + 3.307240000000e-08, + 4.761100000000e-08, + 6.840800000000e-08, + 9.802210000000e-08,  \
+ 1.399280000000e-07, + 1.987290000000e-07, + 2.803210000000e-07, + 3.919410000000e-07, + 5.419990000000e-07,  \
+ 7.396460000000e-07, + 9.940790000000e-07, + 1.313700000000e-06, + 1.705400000000e-06, + 2.174000000000e-06,  \
+ 2.722000000000e-06, + 3.349500000000e-06, + 4.054900000000e-06, + 4.835200000000e-06, + 5.686000000000e-06,  \
+ 6.602500000000e-06, + 7.579800000000e-06, + 8.612700000000e-06, + 9.696300000000e-06, + 1.082580000000e-05,  \
+ 1.199680000000e-05, + 1.320530000000e-05, + 1.444750000000e-05, + 1.572000000000e-05, + 1.701940000000e-05,  \
+ 1.834300000000e-05, + 1.968780000000e-05, + 2.105150000000e-05, + 2.243140000000e-05, + 2.382550000000e-05,  \
+ 2.523150000000e-05, + 2.664750000000e-05, + 2.807140000000e-05, + 2.950160000000e-05, + 3.093610000000e-05,  \
+ 3.237330000000e-05, + 3.381160000000e-05, + 3.524930000000e-05, + 3.668500000000e-05, + 3.811700000000e-05,  \
+ 3.954400000000e-05, + 4.096450000000e-05, + 4.237710000000e-05, + 4.378050000000e-05, + 4.517330000000e-05,  \
+ 4.655430000000e-05, + 4.792220000000e-05, + 4.927570000000e-05, + 5.061360000000e-05, + 5.193470000000e-05,  \
+ 5.323800000000e-05, + 5.452220000000e-05, + 5.578640000000e-05, + 5.702940000000e-05, + 5.825030000000e-05,  \
+ 5.944800000000e-05, + 6.062170000000e-05, + 6.177050000000e-05, + 6.289340000000e-05, + 6.398970000000e-05,  \
+ 6.505860000000e-05, + 6.609950000000e-05, + 6.711160000000e-05, + 6.809430000000e-05, + 6.904710000000e-05 ]

.param id_pred_data_vd0.77=[ \
+ 5.848011652709e-10, + 8.262952477800e-10, + 1.190103436910e-09, + 1.730144287837e-09, + 2.519179780336e-09,  \
+ 3.657423706116e-09, + 5.288180777718e-09, + 7.622086259929e-09, + 1.097103189629e-08, + 1.579298238852e-08,  \
+ 2.275039767241e-08, + 3.278932872774e-08, + 4.724581970095e-08, + 6.799013434033e-08, + 9.760932513814e-08,  \
+ 1.396178367941e-07, + 1.986588620184e-07, + 2.806422043022e-07, + 3.927440809548e-07, + 5.432101278302e-07,  \
+ 7.409346437726e-07, + 9.948558283668e-07, + 1.313259804192e-06, + 1.703123593870e-06, + 2.169599997615e-06,  \
+ 2.715732041452e-06, + 3.342421550769e-06, + 4.048575165143e-06, + 4.831445389755e-06, + 5.686984427484e-06,  \
+ 6.610242480747e-06, + 7.595757124363e-06, + 8.637882801850e-06, + 9.730949095683e-06, + 1.086955030587e-05,  \
+ 1.204867290653e-05, + 1.326360590610e-05, + 1.451015234124e-05, + 1.578452913236e-05, + 1.708344621875e-05,  \
+ 1.840387825723e-05, + 1.974321728994e-05, + 2.109918450515e-05, + 2.246960473713e-05, + 2.385268799117e-05,  \
+ 2.524666248064e-05, + 2.664995110536e-05, + 2.806106360367e-05, + 2.947844528535e-05, + 3.090086640441e-05,  \
+ 3.232683669921e-05, + 3.375500877155e-05, + 3.518397639709e-05, + 3.661242019007e-05, + 3.803895633610e-05,  \
+ 3.946217300836e-05, + 4.088081524969e-05, + 4.229342921462e-05, + 4.369868431240e-05, + 4.509516031248e-05,  \
+ 4.648170870496e-05, + 4.785682242073e-05, + 4.921940337226e-05, + 5.056828063971e-05, + 5.190213203605e-05,  \
+ 5.321992670360e-05, + 5.452072342450e-05, + 5.580337368883e-05, + 5.706714357075e-05, + 5.831118709466e-05,  \
+ 5.953458545264e-05, + 6.073682321585e-05, + 6.191727290570e-05, + 6.307540788839e-05, + 6.421073514502e-05,  \
+ 6.532299696119e-05, + 6.641182357271e-05, + 6.747696286766e-05, + 6.851845966594e-05, + 6.953610107303e-05 ]

* Data table for Id-Vg at Vd = 0.78V
.param vg_data_vd0.78=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.78=[ \
+ 5.828140000000e-10, + 8.426620000000e-10, + 1.218300000000e-09, + 1.761300000000e-09, + 2.546200000000e-09,  \
+ 3.680400000000e-09, + 5.319100000000e-09, + 7.685500000000e-09, + 1.110110000000e-08, + 1.602720000000e-08,  \
+ 2.312350000000e-08, + 3.332940000000e-08, + 4.797380000000e-08, + 6.891810000000e-08, + 9.873590000000e-08,  \
+ 1.409210000000e-07, + 2.000960000000e-07, + 2.821840000000e-07, + 3.944450000000e-07, + 5.453090000000e-07,  \
+ 7.439380000000e-07, + 9.995310000000e-07, + 1.320500000000e-06, + 1.713700000000e-06, + 2.183900000000e-06,  \
+ 2.733500000000e-06, + 3.362700000000e-06, + 4.069900000000e-06, + 4.851900000000e-06, + 5.704500000000e-06,  \
+ 6.622800000000e-06, + 7.601800000000e-06, + 8.636400000000e-06, + 9.721600000000e-06, + 1.085280000000e-05,  \
+ 1.202540000000e-05, + 1.323560000000e-05, + 1.447940000000e-05, + 1.575340000000e-05, + 1.705450000000e-05,  \
+ 1.837970000000e-05, + 1.972610000000e-05, + 2.109140000000e-05, + 2.247300000000e-05, + 2.386870000000e-05,  \
+ 2.527640000000e-05, + 2.669410000000e-05, + 2.811980000000e-05, + 2.955170000000e-05, + 3.098800000000e-05,  \
+ 3.242710000000e-05, + 3.386720000000e-05, + 3.530690000000e-05, + 3.674450000000e-05, + 3.817860000000e-05,  \
+ 3.960770000000e-05, + 4.103030000000e-05, + 4.244520000000e-05, + 4.385090000000e-05, + 4.524610000000e-05,  \
+ 4.662950000000e-05, + 4.799980000000e-05, + 4.935590000000e-05, + 5.069650000000e-05, + 5.202040000000e-05,  \
+ 5.332650000000e-05, + 5.461360000000e-05, + 5.588070000000e-05, + 5.712680000000e-05, + 5.835080000000e-05,  \
+ 5.955180000000e-05, + 6.072870000000e-05, + 6.188080000000e-05, + 6.300720000000e-05, + 6.410690000000e-05,  \
+ 6.517940000000e-05, + 6.622390000000e-05, + 6.723960000000e-05, + 6.822600000000e-05, + 6.918250000000e-05 ]

.param id_pred_data_vd0.78=[ \
+ 5.905694733244e-10, + 8.336247225849e-10, + 1.199641346261e-09, + 1.742952888684e-09, + 2.536929599728e-09,  \
+ 3.682673765937e-09, + 5.324597456280e-09, + 7.674735780228e-09, + 1.104692012532e-08, + 1.590170938925e-08,  \
+ 2.290588827947e-08, + 3.301191938476e-08, + 4.756555256336e-08, + 6.845037816561e-08, + 9.827072489088e-08,  \
+ 1.405601378224e-07, + 1.999811371434e-07, + 2.824589688544e-07, + 3.951783958200e-07, + 5.463805416639e-07,  \
+ 7.449493182321e-07, + 9.997942424889e-07, + 1.319178518315e-06, + 1.710037740850e-06, + 2.177508363275e-06,  \
+ 2.724609794313e-06, + 3.352254152560e-06, + 4.059347002112e-06, + 4.843145425184e-06, + 5.699619996449e-06,  \
+ 6.623836798099e-06, + 7.610347238369e-06, + 8.653459044581e-06, + 9.747567200975e-06, + 1.088721992346e-05,  \
+ 1.206734992593e-05, + 1.328328009549e-05, + 1.453073200537e-05, + 1.580596850545e-05, + 1.710557167826e-05,  \
+ 1.842660742113e-05, + 1.976639417990e-05, + 2.112256253895e-05, + 2.249310771731e-05, + 2.387608736171e-05,  \
+ 2.526976626541e-05, + 2.667268730875e-05, + 2.808323588397e-05, + 2.950002155558e-05, + 3.092168510193e-05,  \
+ 3.234689000237e-05, + 3.377427136002e-05, + 3.520257494529e-05, + 3.663037910883e-05, + 3.805641827057e-05,  \
+ 3.947934455937e-05, + 4.089790374564e-05, + 4.231062310282e-05, + 4.371628245281e-05, + 4.511366445513e-05,  \
+ 4.650127084460e-05, + 4.787792116986e-05, + 4.924246619339e-05, + 5.059366871137e-05, + 5.193036529818e-05,  \
+ 5.325146630639e-05, + 5.455600126879e-05, + 5.584304512013e-05, + 5.711147416150e-05, + 5.836060168804e-05,  \
+ 5.958969559288e-05, + 6.079809187213e-05, + 6.198499031598e-05, + 6.315005608485e-05, + 6.429273300455e-05,  \
+ 6.541265218402e-05, + 6.650944473222e-05, + 6.758298011846e-05, + 6.863298593089e-05, + 6.965943946852e-05 ]

* Data table for Id-Vg at Vd = 0.79V
.param vg_data_vd0.79=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.79=[ \
+ 5.881950000000e-10, + 8.503330000000e-10, + 1.229300000000e-09, + 1.776900000000e-09, + 2.568400000000e-09,  \
+ 3.712000000000e-09, + 5.364000000000e-09, + 7.749500000000e-09, + 1.119200000000e-08, + 1.615620000000e-08,  \
+ 2.330630000000e-08, + 3.358810000000e-08, + 4.833880000000e-08, + 6.943120000000e-08, + 9.945360000000e-08,  \
+ 1.419180000000e-07, + 2.014700000000e-07, + 2.840560000000e-07, + 3.969600000000e-07, + 5.486320000000e-07,  \
+ 7.482450000000e-07, + 1.005000000000e-06, + 1.327300000000e-06, + 1.722000000000e-06, + 2.193700000000e-06,  \
+ 2.745000000000e-06, + 3.375900000000e-06, + 4.084900000000e-06, + 4.868600000000e-06, + 5.722900000000e-06,  \
+ 6.643000000000e-06, + 7.623700000000e-06, + 8.660000000000e-06, + 9.746900000000e-06, + 1.087970000000e-05,  \
+ 1.205400000000e-05, + 1.326570000000e-05, + 1.451120000000e-05, + 1.578680000000e-05, + 1.708950000000e-05,  \
+ 1.841620000000e-05, + 1.976430000000e-05, + 2.113110000000e-05, + 2.251430000000e-05, + 2.391160000000e-05,  \
+ 2.532100000000e-05, + 2.674030000000e-05, + 2.816770000000e-05, + 2.960130000000e-05, + 3.103940000000e-05,  \
+ 3.248030000000e-05, + 3.392230000000e-05, + 3.536390000000e-05, + 3.680340000000e-05, + 3.823950000000e-05,  \
+ 3.967060000000e-05, + 4.109540000000e-05, + 4.251240000000e-05, + 4.392030000000e-05, + 4.531780000000e-05,  \
+ 4.670360000000e-05, + 4.807630000000e-05, + 4.943490000000e-05, + 5.077810000000e-05, + 5.210460000000e-05,  \
+ 5.341340000000e-05, + 5.470340000000e-05, + 5.597340000000e-05, + 5.722240000000e-05, + 5.844940000000e-05,  \
+ 5.965340000000e-05, + 6.083360000000e-05, + 6.198890000000e-05, + 6.311850000000e-05, + 6.422160000000e-05,  \
+ 6.529750000000e-05, + 6.634540000000e-05, + 6.736470000000e-05, + 6.835460000000e-05, + 6.931460000000e-05 ]

.param id_pred_data_vd0.79=[ \
+ 5.964149663029e-10, + 8.410141494331e-10, + 1.209209242736e-09, + 1.755708312068e-09, + 2.554501417062e-09,  \
+ 3.707558926536e-09, + 5.360424792933e-09, + 7.726538839847e-09, + 1.112154780714e-08, + 1.600873702046e-08,  \
+ 2.305917641721e-08, + 3.323157201862e-08, + 4.788158470603e-08, + 6.890583350128e-08, + 9.892544866830e-08,  \
+ 1.414930855503e-07, + 2.012895075154e-07, + 2.842551333515e-07, + 3.975806293965e-07, + 5.495053812865e-07,  \
+ 7.488911086284e-07, + 1.004627417842e-06, + 1.324938942844e-06, + 1.716735191621e-06, + 2.185119585647e-06,  \
+ 2.733109020028e-06, + 3.361595513525e-06, + 4.069505625921e-06, + 4.854108155996e-06, + 5.711372314181e-06,  \
+ 6.636399721174e-06, + 7.623741266798e-06, + 8.667738757140e-06, + 9.762739746293e-06, + 1.090331308660e-05,  \
+ 1.208432293424e-05, + 1.330112561845e-05, + 1.454943600038e-05, + 1.582542303368e-05, + 1.712566234346e-05,  \
+ 1.844717646236e-05, + 1.978730693736e-05, + 2.114372151482e-05, + 2.251424313727e-05, + 2.389706549366e-05,  \
+ 2.529044981202e-05, + 2.669283694559e-05, + 2.810273672367e-05, + 2.951881560875e-05, + 3.093961360719e-05,  \
+ 3.236391788960e-05, + 3.379043802852e-05, + 3.521778013237e-05, + 3.664480322186e-05, + 3.807006167335e-05,  \
+ 3.949248060962e-05, + 4.091061440704e-05, + 4.232320712617e-05, + 4.372903444164e-05, + 4.512673982390e-05,  \
+ 4.651523402572e-05, + 4.789302831341e-05, + 4.925912828185e-05, + 5.061228373961e-05, + 5.195146004553e-05,  \
+ 5.327548460627e-05, + 5.458331128466e-05, + 5.587409512373e-05, + 5.714698541851e-05, + 5.840084406373e-05,  \
+ 5.963516523479e-05, + 6.084918444685e-05, + 6.204222918313e-05, + 6.321379361907e-05, + 6.436345815018e-05,  \
+ 6.549067096785e-05, + 6.659518490778e-05, + 6.767668382963e-05, + 6.873496655317e-05, + 6.976999284234e-05 ]

* Data table for Id-Vg at Vd = 0.80V
.param vg_data_vd0.80=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vd0.80=[ \
+ 5.936180000000e-10, + 8.580630000000e-10, + 1.240300000000e-09, + 1.792600000000e-09, + 2.590800000000e-09,  \
+ 3.743900000000e-09, + 5.409300000000e-09, + 7.813800000000e-09, + 1.128350000000e-08, + 1.628600000000e-08,  \
+ 2.349030000000e-08, + 3.384830000000e-08, + 4.870590000000e-08, + 6.994720000000e-08, + 1.001750000000e-07,  \
+ 1.429210000000e-07, + 2.028520000000e-07, + 2.859370000000e-07, + 3.994860000000e-07, + 5.519670000000e-07,  \
+ 7.525670000000e-07, + 1.010500000000e-06, + 1.334100000000e-06, + 1.730200000000e-06, + 2.203600000000e-06,  \
+ 2.756500000000e-06, + 3.389200000000e-06, + 4.099900000000e-06, + 4.885400000000e-06, + 5.741400000000e-06,  \
+ 6.663200000000e-06, + 7.645600000000e-06, + 8.683600000000e-06, + 9.772200000000e-06, + 1.090660000000e-05,  \
+ 1.208250000000e-05, + 1.329580000000e-05, + 1.454280000000e-05, + 1.582000000000e-05, + 1.712430000000e-05,  \
+ 1.845260000000e-05, + 1.980220000000e-05, + 2.117060000000e-05, + 2.255540000000e-05, + 2.395430000000e-05,  \
+ 2.536530000000e-05, + 2.678630000000e-05, + 2.821530000000e-05, + 2.965070000000e-05, + 3.109050000000e-05,  \
+ 3.253310000000e-05, + 3.397690000000e-05, + 3.542030000000e-05, + 3.686170000000e-05, + 3.829980000000e-05,  \
+ 3.973290000000e-05, + 4.115970000000e-05, + 4.257880000000e-05, + 4.398890000000e-05, + 4.538860000000e-05,  \
+ 4.677660000000e-05, + 4.815180000000e-05, + 4.951280000000e-05, + 5.085840000000e-05, + 5.218750000000e-05,  \
+ 5.349890000000e-05, + 5.479160000000e-05, + 5.606440000000e-05, + 5.731620000000e-05, + 5.854620000000e-05,  \
+ 5.975320000000e-05, + 6.093630000000e-05, + 6.209480000000e-05, + 6.322760000000e-05, + 6.433390000000e-05,  \
+ 6.541310000000e-05, + 6.646430000000e-05, + 6.748690000000e-05, + 6.848020000000e-05, + 6.944370000000e-05 ]

.param id_pred_data_vd0.80=[ \
+ 6.023412879586e-10, + 8.484755120719e-10, + 1.218802214709e-09, + 1.768415280878e-09, + 2.571900559190e-09,  \
+ 3.732099784770e-09, + 5.395648727813e-09, + 7.777414623433e-09, + 1.119488501899e-08, + 1.611405622270e-08,  \
+ 2.321003762518e-08, + 3.344809158534e-08, + 4.819327728001e-08, + 6.935531473573e-08, + 9.957217343981e-08,  \
+ 1.424147171747e-07, + 2.025816684181e-07, + 2.860272616090e-07, + 3.999474756711e-07, + 5.525742380996e-07,  \
+ 7.527518846473e-07, + 1.009341485769e-06, + 1.330529084953e-06, + 1.723200875858e-06, + 2.192418833147e-06,  \
+ 2.741195385170e-06, + 3.370409831405e-06, + 4.079005157109e-06, + 4.864265429205e-06, + 5.722182322643e-06,  \
+ 6.647882401012e-06, + 7.635905785719e-06, + 8.680600149091e-06, + 9.776368824532e-06, + 1.091770172934e-05,  \
+ 1.209952024510e-05, + 1.331709063379e-05, + 1.456612080801e-05, + 1.584275596542e-05, + 1.714355312288e-05,  \
+ 1.846553059295e-05, + 1.980595698114e-05, + 2.116245741490e-05, + 2.253299171571e-05, + 2.391557354713e-05,  \
+ 2.530856290832e-05, + 2.671040128917e-05, + 2.811962040141e-05, + 2.953480579890e-05, + 3.095472056884e-05,  \
+ 3.237798810005e-05, + 3.380342095625e-05, + 3.522973274812e-05, + 3.665566619020e-05, + 3.808014735114e-05,  \
+ 3.950170066673e-05, + 4.091919108760e-05, + 4.233135550749e-05, + 4.373699193820e-05, + 4.513486637734e-05,  \
+ 4.652374482248e-05, + 4.790238454007e-05, + 4.926964757033e-05, + 5.062444251962e-05, + 5.196561687626e-05,  \
+ 5.329204141162e-05, + 5.460293032229e-05, + 5.589705542661e-05, + 5.717368912883e-05, + 5.843203398399e-05,  \
+ 5.967110628262e-05, + 6.089039379731e-05, + 6.208915729076e-05, + 6.326685543172e-05, + 6.442307494581e-05,  \
+ 6.555726868100e-05, + 6.666907574981e-05, + 6.775830406696e-05, + 6.882474990562e-05, + 6.986798834987e-05 ]

* Data table for Id-Vd at Vg = 0.01V
.param vd_data_vg0.01=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.01=[ \
+ 8.817320000000e-11, + 1.486460000000e-10, + 1.899920000000e-10, + 2.183440000000e-10, + 2.383360000000e-10,  \
+ 2.531020000000e-10, + 2.644260000000e-10, + 2.733620000000e-10, + 2.806440000000e-10, + 2.868030000000e-10,  \
+ 2.922060000000e-10, + 2.970960000000e-10, + 3.016350000000e-10, + 3.059300000000e-10, + 3.100540000000e-10,  \
+ 3.140550000000e-10, + 3.179690000000e-10, + 3.218200000000e-10, + 3.256270000000e-10, + 3.294040000000e-10,  \
+ 3.331600000000e-10, + 3.369040000000e-10, + 3.406420000000e-10, + 3.443790000000e-10, + 3.481190000000e-10,  \
+ 3.518670000000e-10, + 3.556230000000e-10, + 3.593920000000e-10, + 3.631750000000e-10, + 3.669740000000e-10,  \
+ 3.707900000000e-10, + 3.746240000000e-10, + 3.784790000000e-10, + 3.823550000000e-10, + 3.862530000000e-10,  \
+ 3.901740000000e-10, + 3.941190000000e-10, + 3.980880000000e-10, + 4.020820000000e-10, + 4.061030000000e-10,  \
+ 4.101500000000e-10, + 4.142250000000e-10, + 4.183270000000e-10, + 4.224580000000e-10, + 4.266170000000e-10,  \
+ 4.308060000000e-10, + 4.350250000000e-10, + 4.392740000000e-10, + 4.435530000000e-10, + 4.478640000000e-10,  \
+ 4.522070000000e-10, + 4.565820000000e-10, + 4.609890000000e-10, + 4.654290000000e-10, + 4.699020000000e-10,  \
+ 4.744090000000e-10, + 4.789500000000e-10, + 4.835250000000e-10, + 4.881350000000e-10, + 4.927800000000e-10,  \
+ 4.974610000000e-10, + 5.021770000000e-10, + 5.069300000000e-10, + 5.117200000000e-10, + 5.165460000000e-10,  \
+ 5.214100000000e-10, + 5.263110000000e-10, + 5.312510000000e-10, + 5.362290000000e-10, + 5.412450000000e-10,  \
+ 5.463010000000e-10, + 5.513960000000e-10, + 5.565310000000e-10, + 5.617060000000e-10, + 5.669220000000e-10,  \
+ 5.721780000000e-10, + 5.774750000000e-10, + 5.828140000000e-10, + 5.881950000000e-10, + 5.936180000000e-10 ]

.param id_pred_data_vg0.01=[ \
+ 8.691662500837e-11, + 1.456778697673e-10, + 1.861711851348e-10, + 2.147539923669e-10, + 2.355277750610e-10,  \
+ 2.511506735914e-10, + 2.633494533555e-10, + 2.732483928014e-10, + 2.815800392852e-10, + 2.888212113916e-10,  \
+ 2.952820987723e-10, + 3.011657589980e-10, + 3.066067399971e-10, + 3.116929470082e-10, + 3.164855377769e-10,  \
+ 3.210287857769e-10, + 3.253566083217e-10, + 3.294980288615e-10, + 3.334754039575e-10, + 3.373139323415e-10,  \
+ 3.410337612308e-10, + 3.446564122989e-10, + 3.482016996958e-10, + 3.516868396503e-10, + 3.551303140448e-10,  \
+ 3.585476271439e-10, + 3.619549160394e-10, + 3.653627578259e-10, + 3.687842653477e-10, + 3.722280150775e-10,  \
+ 3.757040478725e-10, + 3.792177238893e-10, + 3.827742756091e-10, + 3.863791997460e-10, + 3.900331280171e-10,  \
+ 3.937402404119e-10, + 3.975002771384e-10, + 4.013137333558e-10, + 4.051814217476e-10, + 4.091013305896e-10,  \
+ 4.130719388762e-10, + 4.170938128212e-10, + 4.211650606045e-10, + 4.252828578188e-10, + 4.294450794973e-10,  \
+ 4.336522274606e-10, + 4.379006934840e-10, + 4.421913235575e-10, + 4.465209146876e-10, + 4.508873829856e-10,  \
+ 4.552932914015e-10, + 4.597346925372e-10, + 4.642115053466e-10, + 4.687250687585e-10, + 4.732745445546e-10,  \
+ 4.778605822153e-10, + 4.824825555749e-10, + 4.871414427399e-10, + 4.918379326035e-10, + 4.965734157203e-10,  \
+ 5.013510040452e-10, + 5.061688279628e-10, + 5.110306078304e-10, + 5.159360227935e-10, + 5.208905168308e-10,  \
+ 5.258934687724e-10, + 5.309481165838e-10, + 5.360546695421e-10, + 5.412171094621e-10, + 5.464385166576e-10,  \
+ 5.517197532168e-10, + 5.570626759877e-10, + 5.624710763819e-10, + 5.679467607322e-10, + 5.734935026869e-10,  \
+ 5.791107748898e-10, + 5.848011652709e-10, + 5.905694733244e-10, + 5.964149663029e-10, + 6.023412879586e-10 ]

* Data table for Id-Vd at Vg = 0.02V
.param vd_data_vg0.02=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.02=[ \
+ 1.286390000000e-10, + 2.168620000000e-10, + 2.771750000000e-10, + 3.185250000000e-10, + 3.476720000000e-10,  \
+ 3.691890000000e-10, + 3.856790000000e-10, + 3.986810000000e-10, + 4.092660000000e-10, + 4.182090000000e-10,  \
+ 4.260460000000e-10, + 4.331320000000e-10, + 4.397030000000e-10, + 4.459170000000e-10, + 4.518770000000e-10,  \
+ 4.576570000000e-10, + 4.633080000000e-10, + 4.688650000000e-10, + 4.743550000000e-10, + 4.797990000000e-10,  \
+ 4.852120000000e-10, + 4.906050000000e-10, + 4.959880000000e-10, + 5.013680000000e-10, + 5.067510000000e-10,  \
+ 5.121430000000e-10, + 5.175460000000e-10, + 5.229650000000e-10, + 5.284040000000e-10, + 5.338630000000e-10,  \
+ 5.393470000000e-10, + 5.448560000000e-10, + 5.503920000000e-10, + 5.559580000000e-10, + 5.615540000000e-10,  \
+ 5.671820000000e-10, + 5.728430000000e-10, + 5.785380000000e-10, + 5.842690000000e-10, + 5.900360000000e-10,  \
+ 5.958400000000e-10, + 6.016820000000e-10, + 6.075620000000e-10, + 6.134830000000e-10, + 6.194430000000e-10,  \
+ 6.254450000000e-10, + 6.314890000000e-10, + 6.375740000000e-10, + 6.437030000000e-10, + 6.498760000000e-10,  \
+ 6.560930000000e-10, + 6.623550000000e-10, + 6.686620000000e-10, + 6.750150000000e-10, + 6.814150000000e-10,  \
+ 6.878620000000e-10, + 6.943570000000e-10, + 7.008990000000e-10, + 7.074910000000e-10, + 7.141320000000e-10,  \
+ 7.208220000000e-10, + 7.275630000000e-10, + 7.343550000000e-10, + 7.411980000000e-10, + 7.480930000000e-10,  \
+ 7.550400000000e-10, + 7.620400000000e-10, + 7.690930000000e-10, + 7.762000000000e-10, + 7.833610000000e-10,  \
+ 7.905770000000e-10, + 7.978480000000e-10, + 8.051750000000e-10, + 8.125580000000e-10, + 8.199970000000e-10,  \
+ 8.274940000000e-10, + 8.350490000000e-10, + 8.426620000000e-10, + 8.503330000000e-10, + 8.580630000000e-10 ]

.param id_pred_data_vg0.02=[ \
+ 1.277592787119e-10, + 2.137981525152e-10, + 2.727115866463e-10, + 3.139287940712e-10, + 3.435613127323e-10,  \
+ 3.655796465551e-10, + 3.825738437158e-10, + 3.962265537893e-10, + 4.076364046313e-10, + 4.175175760679e-10,  \
+ 4.263325914522e-10, + 4.343790394046e-10, + 4.418489818470e-10, + 4.488720684037e-10, + 4.555236521320e-10,  \
+ 4.618654614319e-10, + 4.679365894766e-10, + 4.737681447153e-10, + 4.793900876265e-10, + 4.848259127499e-10,  \
+ 4.901032779614e-10, + 4.952442411721e-10, + 5.002746061855e-10, + 5.052172546982e-10, + 5.100959099558e-10,  \
+ 5.149317283681e-10, + 5.197448271765e-10, + 5.245532097575e-10, + 5.293776383919e-10, + 5.342262965335e-10,  \
+ 5.391164148438e-10, + 5.440597306006e-10, + 5.490627885685e-10, + 5.541333836234e-10, + 5.592744933836e-10,  \
+ 5.644933320781e-10, + 5.697905169910e-10, + 5.751690634881e-10, + 5.806258840391e-10, + 5.861615193226e-10,  \
+ 5.917750001139e-10, + 5.974638983552e-10, + 6.032243793364e-10, + 6.090571247341e-10, + 6.149545872525e-10,  \
+ 6.209151726111e-10, + 6.269336738640e-10, + 6.330088453410e-10, + 6.391384987925e-10, + 6.453146905727e-10,  \
+ 6.515384731731e-10, + 6.578051348072e-10, + 6.641132033192e-10, + 6.704591681839e-10, + 6.768440197202e-10,  \
+ 6.832605503604e-10, + 6.897126503258e-10, + 6.961959408969e-10, + 7.027135606741e-10, + 7.092601839176e-10,  \
+ 7.158382286931e-10, + 7.224484654955e-10, + 7.290913972557e-10, + 7.357671449881e-10, + 7.424784953525e-10,  \
+ 7.492223574879e-10, + 7.560067527557e-10, + 7.628251985636e-10, + 7.696854420480e-10, + 7.765894149969e-10,  \
+ 7.835373894149e-10, + 7.905324395097e-10, + 7.975775839775e-10, + 8.046725930022e-10, + 8.118217764697e-10,  \
+ 8.190295019972e-10, + 8.262952477800e-10, + 8.336247225849e-10, + 8.410141494331e-10, + 8.484755120719e-10 ]

* Data table for Id-Vd at Vg = 0.03V
.param vd_data_vg0.03=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.03=[ \
+ 1.876680000000e-10, + 3.163730000000e-10, + 4.043540000000e-10, + 4.646600000000e-10, + 5.071520000000e-10,  \
+ 5.385060000000e-10, + 5.625190000000e-10, + 5.814360000000e-10, + 5.968220000000e-10, + 6.098080000000e-10,  \
+ 6.211740000000e-10, + 6.314420000000e-10, + 6.409550000000e-10, + 6.499420000000e-10, + 6.585570000000e-10,  \
+ 6.669050000000e-10, + 6.750620000000e-10, + 6.830790000000e-10, + 6.909970000000e-10, + 6.988440000000e-10,  \
+ 7.066430000000e-10, + 7.144110000000e-10, + 7.221610000000e-10, + 7.299040000000e-10, + 7.376500000000e-10,  \
+ 7.454050000000e-10, + 7.531760000000e-10, + 7.609670000000e-10, + 7.687830000000e-10, + 7.766290000000e-10,  \
+ 7.845060000000e-10, + 7.924190000000e-10, + 8.003700000000e-10, + 8.083600000000e-10, + 8.163930000000e-10,  \
+ 8.244700000000e-10, + 8.325920000000e-10, + 8.407630000000e-10, + 8.489820000000e-10, + 8.572510000000e-10,  \
+ 8.655730000000e-10, + 8.739470000000e-10, + 8.823750000000e-10, + 8.908590000000e-10, + 8.993990000000e-10,  \
+ 9.079960000000e-10, + 9.166520000000e-10, + 9.253670000000e-10, + 9.341420000000e-10, + 9.429780000000e-10,  \
+ 9.518760000000e-10, + 9.608370000000e-10, + 9.698610000000e-10, + 9.789500000000e-10, + 9.881040000000e-10,  \
+ 9.973240000000e-10, + 1.006600000000e-09, + 1.016000000000e-09, + 1.025400000000e-09, + 1.034900000000e-09,  \
+ 1.044400000000e-09, + 1.054100000000e-09, + 1.063800000000e-09, + 1.073500000000e-09, + 1.083400000000e-09,  \
+ 1.093300000000e-09, + 1.103300000000e-09, + 1.113400000000e-09, + 1.123500000000e-09, + 1.133700000000e-09,  \
+ 1.144000000000e-09, + 1.154400000000e-09, + 1.164900000000e-09, + 1.175400000000e-09, + 1.186000000000e-09,  \
+ 1.196700000000e-09, + 1.207500000000e-09, + 1.218300000000e-09, + 1.229300000000e-09, + 1.240300000000e-09 ]

.param id_pred_data_vg0.03=[ \
+ 1.880239075547e-10, + 3.144101157204e-10, + 4.005906539817e-10, + 4.604901349126e-10, + 5.031818961498e-10,  \
+ 5.345861353589e-10, + 5.585687734566e-10, + 5.776620071174e-10, + 5.935148772451e-10, + 6.071995350965e-10,  \
+ 6.194069834820e-10, + 6.305873156975e-10, + 6.410179986815e-10, + 6.508839778263e-10, + 6.602947522083e-10,  \
+ 6.693264964497e-10, + 6.780302364007e-10, + 6.864421031594e-10, + 6.945916841694e-10, + 7.025065418276e-10,  \
+ 7.102143606552e-10, + 7.177449301565e-10, + 7.251252620577e-10, + 7.323830075734e-10, + 7.395511425479e-10,  \
+ 7.466533702427e-10, + 7.537186474948e-10, + 7.607729202164e-10, + 7.678402291766e-10, + 7.749409780544e-10,  \
+ 7.820941472225e-10, + 7.893166298345e-10, + 7.966236270640e-10, + 8.040263832498e-10, + 8.115293437250e-10,  \
+ 8.191473899188e-10, + 8.268767848207e-10, + 8.347267366204e-10, + 8.426942410544e-10, + 8.507754500897e-10,  \
+ 8.589771094414e-10, + 8.672909324048e-10, + 8.757098335366e-10, + 8.842345700089e-10, + 8.928578876244e-10,  \
+ 9.015705559889e-10, + 9.103720000070e-10, + 9.192516614576e-10, + 9.282044133307e-10, + 9.372239651029e-10,  \
+ 9.463009675859e-10, + 9.554319557736e-10, + 9.646088472426e-10, + 9.738298767381e-10, + 9.830831926294e-10,  \
+ 9.923688004676e-10, + 1.001682563562e-09, + 1.011015449137e-09, + 1.020365428817e-09, + 1.029731899749e-09,  \
+ 1.039109743806e-09, + 1.048497166867e-09, + 1.057891874101e-09, + 1.067293169399e-09, + 1.076697897506e-09,  \
+ 1.086110721360e-09, + 1.095523508576e-09, + 1.104942413122e-09, + 1.114367098598e-09, + 1.123796811164e-09,  \
+ 1.133230705941e-09, + 1.142678272004e-09, + 1.152134071480e-09, + 1.161600702293e-09, + 1.171085395324e-09,  \
+ 1.180581779003e-09, + 1.190103436910e-09, + 1.199641346261e-09, + 1.209209242736e-09, + 1.218802214709e-09 ]

* Data table for Id-Vd at Vg = 0.04V
.param vd_data_vg0.04=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.04=[ \
+ 2.737690000000e-10, + 4.615240000000e-10, + 5.898610000000e-10, + 6.778100000000e-10, + 7.397580000000e-10,  \
+ 7.854450000000e-10, + 8.204120000000e-10, + 8.479340000000e-10, + 8.702980000000e-10, + 8.891530000000e-10,  \
+ 9.056390000000e-10, + 9.205150000000e-10, + 9.342860000000e-10, + 9.472830000000e-10, + 9.597330000000e-10,  \
+ 9.717900000000e-10, + 9.835630000000e-10, + 9.951280000000e-10, + 1.006500000000e-09, + 1.017900000000e-09,  \
+ 1.029100000000e-09, + 1.040300000000e-09, + 1.051400000000e-09, + 1.062600000000e-09, + 1.073700000000e-09,  \
+ 1.084900000000e-09, + 1.096000000000e-09, + 1.107200000000e-09, + 1.118500000000e-09, + 1.129700000000e-09,  \
+ 1.141100000000e-09, + 1.152400000000e-09, + 1.163800000000e-09, + 1.175300000000e-09, + 1.186800000000e-09,  \
+ 1.198400000000e-09, + 1.210100000000e-09, + 1.221800000000e-09, + 1.233600000000e-09, + 1.245400000000e-09,  \
+ 1.257400000000e-09, + 1.269400000000e-09, + 1.281400000000e-09, + 1.293600000000e-09, + 1.305800000000e-09,  \
+ 1.318100000000e-09, + 1.330500000000e-09, + 1.343000000000e-09, + 1.355600000000e-09, + 1.368200000000e-09,  \
+ 1.380900000000e-09, + 1.393800000000e-09, + 1.406700000000e-09, + 1.419700000000e-09, + 1.432800000000e-09,  \
+ 1.445900000000e-09, + 1.459200000000e-09, + 1.472600000000e-09, + 1.486100000000e-09, + 1.499600000000e-09,  \
+ 1.513300000000e-09, + 1.527000000000e-09, + 1.540900000000e-09, + 1.554900000000e-09, + 1.568900000000e-09,  \
+ 1.583100000000e-09, + 1.597300000000e-09, + 1.611700000000e-09, + 1.626200000000e-09, + 1.640800000000e-09,  \
+ 1.655500000000e-09, + 1.670200000000e-09, + 1.685200000000e-09, + 1.700200000000e-09, + 1.715300000000e-09,  \
+ 1.730500000000e-09, + 1.745900000000e-09, + 1.761300000000e-09, + 1.776900000000e-09, + 1.792600000000e-09 ]

.param id_pred_data_vg0.04=[ \
+ 2.764217832407e-10, + 4.621736593435e-10, + 5.885365261804e-10, + 6.759600523765e-10, + 7.378449407014e-10,  \
+ 7.829743253751e-10, + 8.171192877882e-10, + 8.440661503073e-10, + 8.662843242746e-10, + 8.853931809938e-10,  \
+ 9.024289759907e-10, + 9.180662630115e-10, + 9.327219041566e-10, + 9.466585915163e-10, + 9.600418460209e-10,  \
+ 9.729694028238e-10, + 9.855070226550e-10, + 9.976935277933e-10, + 1.009561514387e-09, + 1.021143258839e-09,  \
+ 1.032465299922e-09, + 1.043556085989e-09, + 1.054451521654e-09, + 1.065186232552e-09, + 1.075794342498e-09,  \
+ 1.086307985787e-09, + 1.096771313769e-09, + 1.107213698504e-09, + 1.117667665085e-09, + 1.128169158093e-09,  \
+ 1.138734941897e-09, + 1.149402137912e-09, + 1.160186480220e-09, + 1.171101695618e-09, + 1.182167608249e-09,  \
+ 1.193396901300e-09, + 1.204793333986e-09, + 1.216365537182e-09, + 1.228111712326e-09, + 1.240035629735e-09,  \
+ 1.252135515273e-09, + 1.264404061452e-09, + 1.276840879694e-09, + 1.289432924878e-09, + 1.302171770412e-09,  \
+ 1.315056721296e-09, + 1.328069454409e-09, + 1.341199791227e-09, + 1.354440255508e-09, + 1.367773783123e-09,  \
+ 1.381197116679e-09, + 1.394689395084e-09, + 1.408243868184e-09, + 1.421846760330e-09, + 1.435488516943e-09,  \
+ 1.449163384848e-09, + 1.462853558287e-09, + 1.476550872681e-09, + 1.490248864311e-09, + 1.503940172398e-09,  \
+ 1.517610532797e-09, + 1.531256539344e-09, + 1.544870751324e-09, + 1.558451145911e-09, + 1.571988816895e-09,  \
+ 1.585480573496e-09, + 1.598919219248e-09, + 1.612309485921e-09, + 1.625636825153e-09, + 1.638905211543e-09,  \
+ 1.652121233153e-09, + 1.665272080231e-09, + 1.678370409319e-09, + 1.691402609083e-09, + 1.704374308353e-09,  \
+ 1.717290816217e-09, + 1.730144287837e-09, + 1.742952888684e-09, + 1.755708312068e-09, + 1.768415280878e-09 ]

* Data table for Id-Vd at Vg = 0.05V
.param vd_data_vg0.05=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.05=[ \
+ 3.993390000000e-10, + 6.732230000000e-10, + 8.604170000000e-10, + 9.886780000000e-10, + 1.079000000000e-09,  \
+ 1.145600000000e-09, + 1.196500000000e-09, + 1.236500000000e-09, + 1.269000000000e-09, + 1.296400000000e-09,  \
+ 1.320300000000e-09, + 1.341900000000e-09, + 1.361800000000e-09, + 1.380600000000e-09, + 1.398600000000e-09,  \
+ 1.416000000000e-09, + 1.433000000000e-09, + 1.449700000000e-09, + 1.466100000000e-09, + 1.482400000000e-09,  \
+ 1.498600000000e-09, + 1.514700000000e-09, + 1.530700000000e-09, + 1.546800000000e-09, + 1.562800000000e-09,  \
+ 1.578800000000e-09, + 1.594900000000e-09, + 1.611000000000e-09, + 1.627100000000e-09, + 1.643300000000e-09,  \
+ 1.659600000000e-09, + 1.675900000000e-09, + 1.692300000000e-09, + 1.708700000000e-09, + 1.725300000000e-09,  \
+ 1.741900000000e-09, + 1.758600000000e-09, + 1.775400000000e-09, + 1.792300000000e-09, + 1.809300000000e-09,  \
+ 1.826400000000e-09, + 1.843600000000e-09, + 1.860900000000e-09, + 1.878300000000e-09, + 1.895800000000e-09,  \
+ 1.913400000000e-09, + 1.931200000000e-09, + 1.949000000000e-09, + 1.967000000000e-09, + 1.985100000000e-09,  \
+ 2.003300000000e-09, + 2.021600000000e-09, + 2.040100000000e-09, + 2.058700000000e-09, + 2.077400000000e-09,  \
+ 2.096200000000e-09, + 2.115200000000e-09, + 2.134300000000e-09, + 2.153500000000e-09, + 2.172900000000e-09,  \
+ 2.192400000000e-09, + 2.212100000000e-09, + 2.231900000000e-09, + 2.251800000000e-09, + 2.271800000000e-09,  \
+ 2.292100000000e-09, + 2.312400000000e-09, + 2.332900000000e-09, + 2.353600000000e-09, + 2.374400000000e-09,  \
+ 2.395300000000e-09, + 2.416400000000e-09, + 2.437600000000e-09, + 2.459000000000e-09, + 2.480600000000e-09,  \
+ 2.502300000000e-09, + 2.524200000000e-09, + 2.546200000000e-09, + 2.568400000000e-09, + 2.590800000000e-09 ]

.param id_pred_data_vg0.05=[ \
+ 4.053875102272e-10, + 6.780781092175e-10, + 8.634202686153e-10, + 9.912714205029e-10, + 1.081305445183e-09,  \
+ 1.146501560356e-09, + 1.195418430910e-09, + 1.233691904190e-09, + 1.265036475573e-09, + 1.291863949149e-09,  \
+ 1.315746560593e-09, + 1.337685695546e-09, + 1.358314332123e-09, + 1.378021270426e-09, + 1.397039151030e-09,  \
+ 1.415505579416e-09, + 1.433510510296e-09, + 1.451093005755e-09, + 1.468289880791e-09, + 1.485128553469e-09,  \
+ 1.501638053902e-09, + 1.517843903898e-09, + 1.533793603237e-09, + 1.549520618482e-09, + 1.565068519227e-09,  \
+ 1.580484338959e-09, + 1.595814160815e-09, + 1.611109290423e-09, + 1.626417058809e-09, + 1.641777114259e-09,  \
+ 1.657228776430e-09, + 1.672807314890e-09, + 1.688557293988e-09, + 1.704495575794e-09, + 1.720644315917e-09,  \
+ 1.737031478655e-09, + 1.753666230009e-09, + 1.770564566073e-09, + 1.787723742375e-09, + 1.805149807410e-09,  \
+ 1.822843982424e-09, + 1.840802816844e-09, + 1.859015537065e-09, + 1.877474176126e-09, + 1.896167223236e-09,  \
+ 1.915086711435e-09, + 1.934210249743e-09, + 1.953527046794e-09, + 1.973008076916e-09, + 1.992651599281e-09,  \
+ 2.012430089238e-09, + 2.032321031464e-09, + 2.052315135614e-09, + 2.072384583940e-09, + 2.092515205554e-09,  \
+ 2.112682864208e-09, + 2.132868894833e-09, + 2.153061635646e-09, + 2.173242961145e-09, + 2.193393067174e-09,  \
+ 2.213490886138e-09, + 2.233530360662e-09, + 2.253491553361e-09, + 2.273361872085e-09, + 2.293136136533e-09,  \
+ 2.312790639003e-09, + 2.332318453924e-09, + 2.351720462812e-09, + 2.370978913202e-09, + 2.390084574699e-09,  \
+ 2.409027077821e-09, + 2.427813949879e-09, + 2.446434017589e-09, + 2.464884731879e-09, + 2.483153682675e-09,  \
+ 2.501256464171e-09, + 2.519179780336e-09, + 2.536929599728e-09, + 2.554501417062e-09, + 2.571900559190e-09 ]

* Data table for Id-Vd at Vg = 0.06V
.param vd_data_vg0.06=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.06=[ \
+ 5.824360000000e-10, + 9.819230000000e-10, + 1.255000000000e-09, + 1.442000000000e-09, + 1.573700000000e-09,  \
+ 1.670600000000e-09, + 1.744800000000e-09, + 1.803000000000e-09, + 1.850300000000e-09, + 1.890000000000e-09,  \
+ 1.924700000000e-09, + 1.955900000000e-09, + 1.984800000000e-09, + 2.011900000000e-09, + 2.037900000000e-09,  \
+ 2.063100000000e-09, + 2.087600000000e-09, + 2.111600000000e-09, + 2.135300000000e-09, + 2.158800000000e-09,  \
+ 2.182100000000e-09, + 2.205300000000e-09, + 2.228400000000e-09, + 2.251500000000e-09, + 2.274500000000e-09,  \
+ 2.297600000000e-09, + 2.320600000000e-09, + 2.343800000000e-09, + 2.366900000000e-09, + 2.390200000000e-09,  \
+ 2.413500000000e-09, + 2.436900000000e-09, + 2.460400000000e-09, + 2.484000000000e-09, + 2.507800000000e-09,  \
+ 2.531600000000e-09, + 2.555500000000e-09, + 2.579600000000e-09, + 2.603800000000e-09, + 2.628200000000e-09,  \
+ 2.652700000000e-09, + 2.677300000000e-09, + 2.702100000000e-09, + 2.727000000000e-09, + 2.752100000000e-09,  \
+ 2.777300000000e-09, + 2.802700000000e-09, + 2.828200000000e-09, + 2.853900000000e-09, + 2.879800000000e-09,  \
+ 2.905800000000e-09, + 2.932100000000e-09, + 2.958400000000e-09, + 2.985000000000e-09, + 3.011800000000e-09,  \
+ 3.038700000000e-09, + 3.065800000000e-09, + 3.093100000000e-09, + 3.120500000000e-09, + 3.148200000000e-09,  \
+ 3.176000000000e-09, + 3.204100000000e-09, + 3.232300000000e-09, + 3.260800000000e-09, + 3.289400000000e-09,  \
+ 3.318200000000e-09, + 3.347300000000e-09, + 3.376500000000e-09, + 3.405900000000e-09, + 3.435600000000e-09,  \
+ 3.465400000000e-09, + 3.495500000000e-09, + 3.525800000000e-09, + 3.556300000000e-09, + 3.587000000000e-09,  \
+ 3.617900000000e-09, + 3.649100000000e-09, + 3.680400000000e-09, + 3.712000000000e-09, + 3.743900000000e-09 ]

.param id_pred_data_vg0.06=[ \
+ 5.927359936209e-10, + 9.922707278065e-10, + 1.263943296692e-09, + 1.451068811775e-09, + 1.582378850173e-09,  \
+ 1.676932299688e-09, + 1.747377211814e-09, + 1.802077918001e-09, + 1.846566899388e-09, + 1.884461120483e-09,  \
+ 1.918109795440e-09, + 1.949021850578e-09, + 1.978142236680e-09, + 2.006057293613e-09, + 2.033098622789e-09,  \
+ 2.059469892401e-09, + 2.085275978558e-09, + 2.110558767754e-09, + 2.135355146038e-09, + 2.159691447901e-09,  \
+ 2.183587231031e-09, + 2.207068749982e-09, + 2.230175706330e-09, + 2.252957287396e-09, + 2.275459154433e-09,  \
+ 2.297745282931e-09, + 2.319886283075e-09, + 2.341942426654e-09, + 2.363977733566e-09, + 2.386057484927e-09,  \
+ 2.408243142682e-09, + 2.430593895042e-09, + 2.453155838467e-09, + 2.475980522831e-09, + 2.499104811982e-09,  \
+ 2.522554805040e-09, + 2.546367223744e-09, + 2.570560653226e-09, + 2.595146431084e-09, + 2.620133088271e-09,  \
+ 2.645527859002e-09, + 2.671321830405e-09, + 2.697520189443e-09, + 2.724101815232e-09, + 2.751045991012e-09,  \
+ 2.778357330868e-09, + 2.806005010569e-09, + 2.833963463900e-09, + 2.862202781451e-09, + 2.890710115722e-09,  \
+ 2.919458075290e-09, + 2.948404400627e-09, + 2.977524382608e-09, + 3.006796172045e-09, + 3.036177087523e-09,  \
+ 3.065644378353e-09, + 3.095172145251e-09, + 3.124713554570e-09, + 3.154261101201e-09, + 3.183768448878e-09,  \
+ 3.213216577258e-09, + 3.242573010098e-09, + 3.271813979744e-09, + 3.300915238924e-09, + 3.329856057555e-09,  \
+ 3.358607738591e-09, + 3.387153175716e-09, + 3.415466824919e-09, + 3.443535097070e-09, + 3.471336285088e-09,  \
+ 3.498861560480e-09, + 3.526093976802e-09, + 3.553015135438e-09, + 3.579620324601e-09, + 3.605889919989e-09,  \
+ 3.631831315687e-09, + 3.657423706116e-09, + 3.682673765937e-09, + 3.707558926536e-09, + 3.732099784770e-09 ]

* Data table for Id-Vd at Vg = 0.07V
.param vd_data_vg0.07=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.07=[ \
+ 8.493340000000e-10, + 1.432000000000e-09, + 1.830200000000e-09, + 2.102900000000e-09, + 2.294800000000e-09,  \
+ 2.436100000000e-09, + 2.544100000000e-09, + 2.628800000000e-09, + 2.697500000000e-09, + 2.755200000000e-09,  \
+ 2.805400000000e-09, + 2.850700000000e-09, + 2.892400000000e-09, + 2.931700000000e-09, + 2.969200000000e-09,  \
+ 3.005500000000e-09, + 3.040900000000e-09, + 3.075500000000e-09, + 3.109700000000e-09, + 3.143500000000e-09,  \
+ 3.177100000000e-09, + 3.210400000000e-09, + 3.243600000000e-09, + 3.276800000000e-09, + 3.309900000000e-09,  \
+ 3.343100000000e-09, + 3.376200000000e-09, + 3.409400000000e-09, + 3.442700000000e-09, + 3.476100000000e-09,  \
+ 3.509500000000e-09, + 3.543100000000e-09, + 3.576800000000e-09, + 3.610700000000e-09, + 3.644700000000e-09,  \
+ 3.678900000000e-09, + 3.713200000000e-09, + 3.747700000000e-09, + 3.782400000000e-09, + 3.817200000000e-09,  \
+ 3.852300000000e-09, + 3.887600000000e-09, + 3.923000000000e-09, + 3.958700000000e-09, + 3.994600000000e-09,  \
+ 4.030600000000e-09, + 4.067000000000e-09, + 4.103500000000e-09, + 4.140200000000e-09, + 4.177200000000e-09,  \
+ 4.214500000000e-09, + 4.251900000000e-09, + 4.289600000000e-09, + 4.327600000000e-09, + 4.365800000000e-09,  \
+ 4.404200000000e-09, + 4.442900000000e-09, + 4.481900000000e-09, + 4.521100000000e-09, + 4.560600000000e-09,  \
+ 4.600300000000e-09, + 4.640300000000e-09, + 4.680600000000e-09, + 4.721200000000e-09, + 4.762000000000e-09,  \
+ 4.803100000000e-09, + 4.844500000000e-09, + 4.886200000000e-09, + 4.928100000000e-09, + 4.970400000000e-09,  \
+ 5.012900000000e-09, + 5.055800000000e-09, + 5.098900000000e-09, + 5.142300000000e-09, + 5.186000000000e-09,  \
+ 5.230100000000e-09, + 5.274400000000e-09, + 5.319100000000e-09, + 5.364000000000e-09, + 5.409300000000e-09 ]

.param id_pred_data_vg0.07=[ \
+ 8.640822102279e-10, + 1.448235451562e-09, + 1.846051844723e-09, + 2.120021065366e-09, + 2.311887747908e-09,  \
+ 2.449504279411e-09, + 2.551454514332e-09, + 2.630122253322e-09, + 2.693707017443e-09, + 2.747617777743e-09,  \
+ 2.795372129327e-09, + 2.839225174966e-09, + 2.880601872590e-09, + 2.920371890980e-09, + 2.959027156635e-09,  \
+ 2.996842454195e-09, + 3.033966198274e-09, + 3.070429031027e-09, + 3.106259782726e-09, + 3.141463622569e-09,  \
+ 3.176034368835e-09, + 3.210004457799e-09, + 3.243395347852e-09, + 3.276252016349e-09, + 3.308640028621e-09,  \
+ 3.340643726091e-09, + 3.372351358166e-09, + 3.403836110749e-09, + 3.435200834900e-09, + 3.466552112030e-09,  \
+ 3.497969913724e-09, + 3.529545722358e-09, + 3.561350681025e-09, + 3.593485633502e-09, + 3.625995015355e-09,  \
+ 3.658965290754e-09, + 3.692413317324e-09, + 3.726386825775e-09, + 3.760922133722e-09, + 3.796047209903e-09,  \
+ 3.831764763262e-09, + 3.868083933156e-09, + 3.905006042970e-09, + 3.942523818523e-09, + 3.980623430877e-09,  \
+ 4.019290678059e-09, + 4.058489366798e-09, + 4.098192505353e-09, + 4.138382188046e-09, + 4.179002033311e-09,  \
+ 4.220022731261e-09, + 4.261425061713e-09, + 4.303135741068e-09, + 4.345124580141e-09, + 4.387348750967e-09,  \
+ 4.429760522839e-09, + 4.472307750802e-09, + 4.514941576161e-09, + 4.557643737968e-09, + 4.600340908212e-09,  \
+ 4.642998128190e-09, + 4.685568750773e-09, + 4.728011901989e-09, + 4.770283794642e-09, + 4.812355269834e-09,  \
+ 4.854167041657e-09, + 4.895694094564e-09, + 4.936890700691e-09, + 4.977737262379e-09, + 5.018193105499e-09,  \
+ 5.058234582300e-09, + 5.097817528110e-09, + 5.136934695393e-09, + 5.175548531966e-09, + 5.213639520107e-09,  \
+ 5.251187324973e-09, + 5.288180777718e-09, + 5.324597456280e-09, + 5.360424792933e-09, + 5.395648727813e-09 ]

* Data table for Id-Vd at Vg = 0.08V
.param vd_data_vg0.08=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.08=[ \
+ 1.238200000000e-09, + 2.087800000000e-09, + 2.668500000000e-09, + 3.066100000000e-09, + 3.345900000000e-09,  \
+ 3.551800000000e-09, + 3.708900000000e-09, + 3.832200000000e-09, + 3.931900000000e-09, + 4.015700000000e-09,  \
+ 4.088600000000e-09, + 4.154000000000e-09, + 4.214400000000e-09, + 4.271200000000e-09, + 4.325400000000e-09,  \
+ 4.377800000000e-09, + 4.428800000000e-09, + 4.478700000000e-09, + 4.528000000000e-09, + 4.576600000000e-09,  \
+ 4.624900000000e-09, + 4.672900000000e-09, + 4.720600000000e-09, + 4.768300000000e-09, + 4.815900000000e-09,  \
+ 4.863500000000e-09, + 4.911100000000e-09, + 4.958800000000e-09, + 5.006500000000e-09, + 5.054400000000e-09,  \
+ 5.102400000000e-09, + 5.150600000000e-09, + 5.198900000000e-09, + 5.247400000000e-09, + 5.296200000000e-09,  \
+ 5.345100000000e-09, + 5.394300000000e-09, + 5.443700000000e-09, + 5.493300000000e-09, + 5.543300000000e-09,  \
+ 5.593400000000e-09, + 5.643900000000e-09, + 5.694600000000e-09, + 5.745600000000e-09, + 5.796900000000e-09,  \
+ 5.848500000000e-09, + 5.900400000000e-09, + 5.952700000000e-09, + 6.005200000000e-09, + 6.058000000000e-09,  \
+ 6.111200000000e-09, + 6.164700000000e-09, + 6.218600000000e-09, + 6.272800000000e-09, + 6.327300000000e-09,  \
+ 6.382200000000e-09, + 6.437400000000e-09, + 6.493000000000e-09, + 6.548900000000e-09, + 6.605200000000e-09,  \
+ 6.661900000000e-09, + 6.719000000000e-09, + 6.776400000000e-09, + 6.834200000000e-09, + 6.892400000000e-09,  \
+ 6.951000000000e-09, + 7.010000000000e-09, + 7.069300000000e-09, + 7.129100000000e-09, + 7.189300000000e-09,  \
+ 7.249800000000e-09, + 7.310800000000e-09, + 7.372200000000e-09, + 7.434000000000e-09, + 7.496300000000e-09,  \
+ 7.558900000000e-09, + 7.622000000000e-09, + 7.685500000000e-09, + 7.749500000000e-09, + 7.813800000000e-09 ]

.param id_pred_data_vg0.08=[ \
+ 1.256348838297e-09, + 2.108810548407e-09, + 2.690773897029e-09, + 3.091963662882e-09, + 3.372719703520e-09,  \
+ 3.573605624752e-09, + 3.721830488246e-09, + 3.835617974346e-09, + 3.927132858905e-09, + 4.004414932979e-09,  \
+ 4.072723029935e-09, + 4.135463171906e-09, + 4.194753842057e-09, + 4.251896967844e-09, + 4.307617729182e-09,  \
+ 4.362318293261e-09, + 4.416163097432e-09, + 4.469186620781e-09, + 4.521391847589e-09, + 4.572720868623e-09,  \
+ 4.623148051053e-09, + 4.672640940839e-09, + 4.721210125069e-09, + 4.768891841422e-09, + 4.815769116817e-09,  \
+ 4.861896485409e-09, + 4.907406641053e-09, + 4.952429222271e-09, + 4.997072604596e-09, + 5.041504813619e-09,  \
+ 5.085828647111e-09, + 5.130231102157e-09, + 5.174801387398e-09, + 5.219682002178e-09, + 5.264995195375e-09,  \
+ 5.310821862281e-09, + 5.357264916128e-09, + 5.404401353104e-09, + 5.452283584617e-09, + 5.500958977223e-09,  \
+ 5.550462764958e-09, + 5.600850236931e-09, + 5.652090955266e-09, + 5.704239569582e-09, + 5.757222298897e-09,  \
+ 5.811073968687e-09, + 5.865755774437e-09, + 5.921230012973e-09, + 5.977461272622e-09, + 6.034417410206e-09,  \
+ 6.092035889083e-09, + 6.150278686334e-09, + 6.209067962004e-09, + 6.268362628958e-09, + 6.328081481044e-09,  \
+ 6.388182001160e-09, + 6.448579776830e-09, + 6.509221179840e-09, + 6.570033344033e-09, + 6.630962978704e-09,  \
+ 6.691913476686e-09, + 6.752845180813e-09, + 6.813663473437e-09, + 6.874320206407e-09, + 6.934776042300e-09,  \
+ 6.994934871329e-09, + 7.054749486812e-09, + 7.114141382658e-09, + 7.173084073386e-09, + 7.231520360307e-09,  \
+ 7.289389429843e-09, + 7.346628265736e-09, + 7.403199102640e-09, + 7.459089541584e-09, + 7.514216582294e-09,  \
+ 7.568549627024e-09, + 7.622086259929e-09, + 7.674735780228e-09, + 7.726538839847e-09, + 7.777414623433e-09 ]

* Data table for Id-Vd at Vg = 0.09V
.param vd_data_vg0.09=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.09=[ \
+ 1.804500000000e-09, + 3.043000000000e-09, + 3.889600000000e-09, + 4.469400000000e-09, + 4.877100000000e-09,  \
+ 5.177000000000e-09, + 5.405800000000e-09, + 5.585100000000e-09, + 5.730000000000e-09, + 5.851500000000e-09,  \
+ 5.957200000000e-09, + 6.052000000000e-09, + 6.139300000000e-09, + 6.221300000000e-09, + 6.299600000000e-09,  \
+ 6.375100000000e-09, + 6.448600000000e-09, + 6.520600000000e-09, + 6.591500000000e-09, + 6.661500000000e-09,  \
+ 6.730900000000e-09, + 6.799900000000e-09, + 6.868600000000e-09, + 6.937000000000e-09, + 7.005400000000e-09,  \
+ 7.073700000000e-09, + 7.142000000000e-09, + 7.210400000000e-09, + 7.278900000000e-09, + 7.347500000000e-09,  \
+ 7.416400000000e-09, + 7.485400000000e-09, + 7.554600000000e-09, + 7.624200000000e-09, + 7.693900000000e-09,  \
+ 7.764000000000e-09, + 7.834400000000e-09, + 7.905100000000e-09, + 7.976200000000e-09, + 8.047600000000e-09,  \
+ 8.119400000000e-09, + 8.191500000000e-09, + 8.264000000000e-09, + 8.336900000000e-09, + 8.410300000000e-09,  \
+ 8.484000000000e-09, + 8.558200000000e-09, + 8.632800000000e-09, + 8.707800000000e-09, + 8.783200000000e-09,  \
+ 8.859200000000e-09, + 8.935500000000e-09, + 9.012400000000e-09, + 9.089700000000e-09, + 9.167500000000e-09,  \
+ 9.245700000000e-09, + 9.324500000000e-09, + 9.403800000000e-09, + 9.483500000000e-09, + 9.563800000000e-09,  \
+ 9.644600000000e-09, + 9.725900000000e-09, + 9.807700000000e-09, + 9.890000000000e-09, + 9.972900000000e-09,  \
+ 1.005630000000e-08, + 1.014030000000e-08, + 1.022480000000e-08, + 1.030980000000e-08, + 1.039550000000e-08,  \
+ 1.048170000000e-08, + 1.056840000000e-08, + 1.065570000000e-08, + 1.074360000000e-08, + 1.083210000000e-08,  \
+ 1.092120000000e-08, + 1.101090000000e-08, + 1.110110000000e-08, + 1.119200000000e-08, + 1.128350000000e-08 ]

.param id_pred_data_vg0.09=[ \
+ 1.822785691274e-09, + 3.064841394007e-09, + 3.915456119330e-09, + 4.502927026806e-09, + 4.914190654404e-09,  \
+ 5.208061821804e-09, + 5.424245301811e-09, + 5.589569127551e-09, + 5.721949634108e-09, + 5.833383909248e-09,  \
+ 5.931702666828e-09, + 6.022046221688e-09, + 6.107592867011e-09, + 6.190274035589e-09, + 6.271229935351e-09,  \
+ 6.350998660309e-09, + 6.429819379150e-09, + 6.507665446520e-09, + 6.584486236250e-09, + 6.660125961844e-09,  \
+ 6.734497439709e-09, + 6.807462966663e-09, + 6.878983320746e-09, + 6.949053812377e-09, + 7.017709968693e-09,  \
+ 7.085022986075e-09, + 7.151138241568e-09, + 7.216222570605e-09, + 7.280425489142e-09, + 7.343969699036e-09,  \
+ 7.407039124274e-09, + 7.469853926523e-09, + 7.532623591544e-09, + 7.595519697645e-09, + 7.658769707319e-09,  \
+ 7.722529815624e-09, + 7.786928168940e-09, + 7.852147305698e-09, + 7.918256663686e-09, + 7.985381955677e-09,  \
+ 8.053632960525e-09, + 8.123009571648e-09, + 8.193588616479e-09, + 8.265401660879e-09, + 8.338450729894e-09,  \
+ 8.412739234132e-09, + 8.488243281590e-09, + 8.564940117139e-09, + 8.642782525214e-09, + 8.721740663020e-09,  \
+ 8.801760920107e-09, + 8.882741511229e-09, + 8.964639821585e-09, + 9.047367655057e-09, + 9.130843903193e-09,  \
+ 9.214979570515e-09, + 9.299709482491e-09, + 9.384888102204e-09, + 9.470488571139e-09, + 9.556348246065e-09,  \
+ 9.642403373533e-09, + 9.728549166255e-09, + 9.814745016712e-09, + 9.900795703288e-09, + 9.986686499985e-09,  \
+ 1.007228316752e-08, + 1.015752099320e-08, + 1.024229263180e-08, + 1.032648361488e-08, + 1.041009198843e-08,  \
+ 1.049295711653e-08, + 1.057502885260e-08, + 1.065625546914e-08, + 1.073650111039e-08, + 1.081578759887e-08,  \
+ 1.089397212439e-08, + 1.097103189629e-08, + 1.104692012532e-08, + 1.112154780714e-08, + 1.119488501899e-08 ]

* Data table for Id-Vd at Vg = 0.10V
.param vd_data_vg0.10=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.10=[ \
+ 2.628400000000e-09, + 4.433200000000e-09, + 5.667200000000e-09, + 6.512300000000e-09, + 7.106500000000e-09,  \
+ 7.543300000000e-09, + 7.876200000000e-09, + 8.137000000000e-09, + 8.347500000000e-09, + 8.523800000000e-09,  \
+ 8.676900000000e-09, + 8.814100000000e-09, + 8.940300000000e-09, + 9.058800000000e-09, + 9.171700000000e-09,  \
+ 9.280600000000e-09, + 9.386500000000e-09, + 9.490100000000e-09, + 9.592100000000e-09, + 9.692800000000e-09,  \
+ 9.792600000000e-09, + 9.891700000000e-09, + 9.990300000000e-09, + 1.008860000000e-08, + 1.018670000000e-08,  \
+ 1.028470000000e-08, + 1.038270000000e-08, + 1.048070000000e-08, + 1.057890000000e-08, + 1.067720000000e-08,  \
+ 1.077580000000e-08, + 1.087470000000e-08, + 1.097380000000e-08, + 1.107330000000e-08, + 1.117320000000e-08,  \
+ 1.127340000000e-08, + 1.137410000000e-08, + 1.147530000000e-08, + 1.157680000000e-08, + 1.167890000000e-08,  \
+ 1.178150000000e-08, + 1.188450000000e-08, + 1.198810000000e-08, + 1.209230000000e-08, + 1.219700000000e-08,  \
+ 1.230220000000e-08, + 1.240810000000e-08, + 1.251450000000e-08, + 1.262160000000e-08, + 1.272920000000e-08,  \
+ 1.283750000000e-08, + 1.294640000000e-08, + 1.305600000000e-08, + 1.316620000000e-08, + 1.327700000000e-08,  \
+ 1.338860000000e-08, + 1.350080000000e-08, + 1.361370000000e-08, + 1.372730000000e-08, + 1.384160000000e-08,  \
+ 1.395660000000e-08, + 1.407230000000e-08, + 1.418870000000e-08, + 1.430590000000e-08, + 1.442380000000e-08,  \
+ 1.454250000000e-08, + 1.466190000000e-08, + 1.478210000000e-08, + 1.490300000000e-08, + 1.502480000000e-08,  \
+ 1.514730000000e-08, + 1.527060000000e-08, + 1.539460000000e-08, + 1.551950000000e-08, + 1.564520000000e-08,  \
+ 1.577170000000e-08, + 1.589900000000e-08, + 1.602720000000e-08, + 1.615620000000e-08, + 1.628600000000e-08 ]

.param id_pred_data_vg0.10=[ \
+ 2.640145453370e-09, + 4.447545052244e-09, + 5.689836655165e-09, + 6.549920499310e-09, + 7.152573999747e-09,  \
+ 7.582889622881e-09, + 7.898721321453e-09, + 8.139339229274e-09, + 8.331265277661e-09, + 8.492235537005e-09,  \
+ 8.634034074362e-09, + 8.764331766997e-09, + 8.887953057979e-09, + 9.007895442892e-09, + 9.125821165412e-09,  \
+ 9.242517080565e-09, + 9.358365637979e-09, + 9.473222206680e-09, + 9.586969795805e-09, + 9.699265035579e-09,  \
+ 9.809836996055e-09, + 9.918449634938e-09, + 1.002491046620e-08, + 1.012907347331e-08, + 1.023094320374e-08,  \
+ 1.033057422717e-08, + 1.042803059903e-08, + 1.052352047282e-08, + 1.061722979756e-08, + 1.070948876247e-08,  \
+ 1.080051323044e-08, + 1.089065335691e-08, + 1.098015694367e-08, + 1.106938988471e-08, + 1.115860897016e-08,  \
+ 1.124811475961e-08, + 1.133812858711e-08, + 1.142892536166e-08, + 1.152068755061e-08, + 1.161361069535e-08,  \
+ 1.170786905647e-08, + 1.180356772323e-08, + 1.190079082392e-08, + 1.199964785314e-08, + 1.210018245601e-08,  \
+ 1.220242047850e-08, + 1.230632506122e-08, + 1.241198077651e-08, + 1.251931694313e-08, + 1.262824600445e-08,  \
+ 1.273876103269e-08, + 1.285074226587e-08, + 1.296412964535e-08, + 1.307885096224e-08, + 1.319474192130e-08,  \
+ 1.331172782670e-08, + 1.342971851059e-08, + 1.354853942814e-08, + 1.366807559577e-08, + 1.378820257969e-08,  \
+ 1.390881058327e-08, + 1.402975367881e-08, + 1.415087327317e-08, + 1.427200118087e-08, + 1.439306798190e-08,  \
+ 1.451393991658e-08, + 1.463442101723e-08, + 1.475447199084e-08, + 1.487387999433e-08, + 1.499253396986e-08,  \
+ 1.511037650559e-08, + 1.522722811842e-08, + 1.534295959615e-08, + 1.545749512388e-08, + 1.557075401948e-08,  \
+ 1.568259285989e-08, + 1.579298238852e-08, + 1.590170938925e-08, + 1.600873702046e-08, + 1.611405622270e-08 ]

* Data table for Id-Vd at Vg = 0.11V
.param vd_data_vg0.11=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.11=[ \
+ 3.825400000000e-09, + 6.454000000000e-09, + 8.252200000000e-09, + 9.483700000000e-09, + 1.034930000000e-08,  \
+ 1.098530000000e-08, + 1.146990000000e-08, + 1.184890000000e-08, + 1.215470000000e-08, + 1.241040000000e-08,  \
+ 1.263210000000e-08, + 1.283060000000e-08, + 1.301300000000e-08, + 1.318400000000e-08, + 1.334680000000e-08,  \
+ 1.350370000000e-08, + 1.365610000000e-08, + 1.380520000000e-08, + 1.395180000000e-08, + 1.409650000000e-08,  \
+ 1.423980000000e-08, + 1.438210000000e-08, + 1.452360000000e-08, + 1.466460000000e-08, + 1.480520000000e-08,  \
+ 1.494560000000e-08, + 1.508600000000e-08, + 1.522640000000e-08, + 1.536700000000e-08, + 1.550780000000e-08,  \
+ 1.564880000000e-08, + 1.579020000000e-08, + 1.593200000000e-08, + 1.607430000000e-08, + 1.621710000000e-08,  \
+ 1.636030000000e-08, + 1.650420000000e-08, + 1.664860000000e-08, + 1.679370000000e-08, + 1.693940000000e-08,  \
+ 1.708580000000e-08, + 1.723290000000e-08, + 1.738080000000e-08, + 1.752930000000e-08, + 1.767860000000e-08,  \
+ 1.782870000000e-08, + 1.797960000000e-08, + 1.813140000000e-08, + 1.828390000000e-08, + 1.843730000000e-08,  \
+ 1.859150000000e-08, + 1.874670000000e-08, + 1.890270000000e-08, + 1.905960000000e-08, + 1.921740000000e-08,  \
+ 1.937610000000e-08, + 1.953580000000e-08, + 1.969640000000e-08, + 1.985800000000e-08, + 2.002050000000e-08,  \
+ 2.018400000000e-08, + 2.034850000000e-08, + 2.051410000000e-08, + 2.068060000000e-08, + 2.084810000000e-08,  \
+ 2.101670000000e-08, + 2.118630000000e-08, + 2.135700000000e-08, + 2.152870000000e-08, + 2.170150000000e-08,  \
+ 2.187540000000e-08, + 2.205030000000e-08, + 2.222640000000e-08, + 2.240360000000e-08, + 2.258180000000e-08,  \
+ 2.276120000000e-08, + 2.294180000000e-08, + 2.312350000000e-08, + 2.330630000000e-08, + 2.349030000000e-08 ]

.param id_pred_data_vg0.11=[ \
+ 3.818819322987e-09, + 6.446107931879e-09, + 8.259114565590e-09, + 9.517726198283e-09, + 1.040068298153e-08,  \
+ 1.103074623643e-08, + 1.149206738660e-08, + 1.184209281746e-08, + 1.211989740568e-08, + 1.235191149362e-08,  \
+ 1.255567831038e-08, + 1.274283675912e-08, + 1.292070187731e-08, + 1.309384259685e-08, + 1.326480365549e-08,  \
+ 1.343486133010e-08, + 1.360450426091e-08, + 1.377352248255e-08, + 1.394167092883e-08, + 1.410836460991e-08,  \
+ 1.427298364831e-08, + 1.443505723842e-08, + 1.459417227068e-08, + 1.474992075146e-08, + 1.490224121881e-08,  \
+ 1.505092207310e-08, + 1.519606648515e-08, + 1.533779297347e-08, + 1.547640827937e-08, + 1.561214304502e-08,  \
+ 1.574537680682e-08, + 1.587660335645e-08, + 1.600616844399e-08, + 1.613452361937e-08, + 1.626217951411e-08,  \
+ 1.638946386606e-08, + 1.651684080173e-08, + 1.664472904395e-08, + 1.677343895778e-08, + 1.690331288273e-08,  \
+ 1.703458920588e-08, + 1.716750645642e-08, + 1.730227719321e-08, + 1.743914879171e-08, + 1.757807979175e-08,  \
+ 1.771930115524e-08, + 1.786282172844e-08, + 1.800865845780e-08, + 1.815680853667e-08, + 1.830724372098e-08,  \
+ 1.845999214822e-08, + 1.861480811272e-08, + 1.877178529952e-08, + 1.893071235770e-08, + 1.909142728351e-08,  \
+ 1.925397242530e-08, + 1.941796515581e-08, + 1.958337939811e-08, + 1.975001975296e-08, + 1.991767177856e-08,  \
+ 2.008626413641e-08, + 2.025555090768e-08, + 2.042527651014e-08, + 2.059531880150e-08, + 2.076550824626e-08,  \
+ 2.093558158833e-08, + 2.110550518353e-08, + 2.127490731141e-08, + 2.144364760426e-08, + 2.161166214876e-08,  \
+ 2.177862214126e-08, + 2.194444562065e-08, + 2.210895338806e-08, + 2.227195778914e-08, + 2.243330587959e-08,  \
+ 2.259284229922e-08, + 2.275039767241e-08, + 2.290588827947e-08, + 2.305917641721e-08, + 2.321003762518e-08 ]

* Data table for Id-Vd at Vg = 0.12V
.param vd_data_vg0.12=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.12=[ \
+ 5.561200000000e-09, + 9.386900000000e-09, + 1.200550000000e-08, + 1.379950000000e-08, + 1.506010000000e-08,  \
+ 1.598600000000e-08, + 1.669080000000e-08, + 1.724170000000e-08, + 1.768560000000e-08, + 1.805630000000e-08,  \
+ 1.837730000000e-08, + 1.866420000000e-08, + 1.892760000000e-08, + 1.917420000000e-08, + 1.940880000000e-08,  \
+ 1.963450000000e-08, + 1.985370000000e-08, + 2.006800000000e-08, + 2.027850000000e-08, + 2.048620000000e-08,  \
+ 2.069180000000e-08, + 2.089580000000e-08, + 2.109860000000e-08, + 2.130050000000e-08, + 2.150190000000e-08,  \
+ 2.170290000000e-08, + 2.190370000000e-08, + 2.210450000000e-08, + 2.230550000000e-08, + 2.250670000000e-08,  \
+ 2.270830000000e-08, + 2.291030000000e-08, + 2.311290000000e-08, + 2.331600000000e-08, + 2.351970000000e-08,  \
+ 2.372420000000e-08, + 2.392940000000e-08, + 2.413540000000e-08, + 2.434230000000e-08, + 2.455000000000e-08,  \
+ 2.475870000000e-08, + 2.496830000000e-08, + 2.517890000000e-08, + 2.539050000000e-08, + 2.560310000000e-08,  \
+ 2.581680000000e-08, + 2.603160000000e-08, + 2.624750000000e-08, + 2.646450000000e-08, + 2.668270000000e-08,  \
+ 2.690200000000e-08, + 2.712260000000e-08, + 2.734440000000e-08, + 2.756740000000e-08, + 2.779160000000e-08,  \
+ 2.801710000000e-08, + 2.824390000000e-08, + 2.847210000000e-08, + 2.870150000000e-08, + 2.893220000000e-08,  \
+ 2.916430000000e-08, + 2.939780000000e-08, + 2.963260000000e-08, + 2.986890000000e-08, + 3.010650000000e-08,  \
+ 3.034550000000e-08, + 3.058600000000e-08, + 3.082790000000e-08, + 3.107130000000e-08, + 3.131620000000e-08,  \
+ 3.156250000000e-08, + 3.181030000000e-08, + 3.205970000000e-08, + 3.231050000000e-08, + 3.256290000000e-08,  \
+ 3.281690000000e-08, + 3.307240000000e-08, + 3.332940000000e-08, + 3.358810000000e-08, + 3.384830000000e-08 ]

.param id_pred_data_vg0.12=[ \
+ 5.517154022527e-09, + 9.332759987046e-09, + 1.197685151055e-08, + 1.381769607178e-08, + 1.511071019422e-08,  \
+ 1.603267492101e-08, + 1.670562255640e-08, + 1.721363787510e-08, + 1.761427739666e-08, + 1.794673067934e-08,  \
+ 1.823736724305e-08, + 1.850365833889e-08, + 1.875687033248e-08, + 1.900403105992e-08, + 1.924907380157e-08,  \
+ 1.949415946001e-08, + 1.973997584059e-08, + 1.998634346023e-08, + 2.023265295747e-08, + 2.047804059657e-08,  \
+ 2.072140880216e-08, + 2.096198315371e-08, + 2.119878573126e-08, + 2.143110521047e-08, + 2.165849366520e-08,  \
+ 2.188059127661e-08, + 2.209728720004e-08, + 2.230856949836e-08, + 2.251464884750e-08, + 2.271587931091e-08,  \
+ 2.291266660848e-08, + 2.310552190465e-08, + 2.329505804255e-08, + 2.348186171730e-08, + 2.366656737252e-08,  \
+ 2.384980405168e-08, + 2.403232059578e-08, + 2.421456457569e-08, + 2.439711067836e-08, + 2.458057508647e-08,  \
+ 2.476523725647e-08, + 2.495176673278e-08, + 2.514030821743e-08, + 2.533125893933e-08, + 2.552478548523e-08,  \
+ 2.572121488242e-08, + 2.592064699769e-08, + 2.612314972339e-08, + 2.632886200615e-08, + 2.653769293204e-08,  \
+ 2.674962043869e-08, + 2.696469991292e-08, + 2.718275560198e-08, + 2.740379507316e-08, + 2.762743189777e-08,  \
+ 2.785367115621e-08, + 2.808239518259e-08, + 2.831324607655e-08, + 2.854600186453e-08, + 2.878063654066e-08,  \
+ 2.901671905420e-08, + 2.925407272869e-08, + 2.949239124916e-08, + 2.973145228680e-08, + 2.997107930724e-08,  \
+ 3.021090194011e-08, + 3.045064620011e-08, + 3.069014013590e-08, + 3.092901508239e-08, + 3.116706643880e-08,  \
+ 3.140407383029e-08, + 3.163968415265e-08, + 3.187371014235e-08, + 3.210601505543e-08, + 3.233607781539e-08,  \
+ 3.256398912299e-08, + 3.278932872774e-08, + 3.301191938476e-08, + 3.323157201862e-08, + 3.344809158534e-08 ]

* Data table for Id-Vd at Vg = 0.13V
.param vd_data_vg0.13=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.13=[ \
+ 8.071600000000e-09, + 1.363300000000e-08, + 1.744360000000e-08, + 2.005540000000e-08, + 2.189060000000e-08,  \
+ 2.323780000000e-08, + 2.426260000000e-08, + 2.506280000000e-08, + 2.570680000000e-08, + 2.624390000000e-08,  \
+ 2.670820000000e-08, + 2.712270000000e-08, + 2.750250000000e-08, + 2.785770000000e-08, + 2.819520000000e-08,  \
+ 2.851970000000e-08, + 2.883450000000e-08, + 2.914200000000e-08, + 2.944390000000e-08, + 2.974150000000e-08,  \
+ 3.003590000000e-08, + 3.032790000000e-08, + 3.061800000000e-08, + 3.090670000000e-08, + 3.119450000000e-08,  \
+ 3.148170000000e-08, + 3.176860000000e-08, + 3.205530000000e-08, + 3.234210000000e-08, + 3.262920000000e-08,  \
+ 3.291670000000e-08, + 3.320470000000e-08, + 3.349340000000e-08, + 3.378280000000e-08, + 3.407300000000e-08,  \
+ 3.436420000000e-08, + 3.465640000000e-08, + 3.494960000000e-08, + 3.524390000000e-08, + 3.553950000000e-08,  \
+ 3.583620000000e-08, + 3.613430000000e-08, + 3.643360000000e-08, + 3.673430000000e-08, + 3.703640000000e-08,  \
+ 3.734000000000e-08, + 3.764500000000e-08, + 3.795160000000e-08, + 3.825970000000e-08, + 3.856930000000e-08,  \
+ 3.888060000000e-08, + 3.919350000000e-08, + 3.950800000000e-08, + 3.982430000000e-08, + 4.014220000000e-08,  \
+ 4.046190000000e-08, + 4.078330000000e-08, + 4.110650000000e-08, + 4.143140000000e-08, + 4.175820000000e-08,  \
+ 4.208690000000e-08, + 4.241740000000e-08, + 4.274980000000e-08, + 4.308410000000e-08, + 4.342030000000e-08,  \
+ 4.375840000000e-08, + 4.409850000000e-08, + 4.444060000000e-08, + 4.478460000000e-08, + 4.513070000000e-08,  \
+ 4.547880000000e-08, + 4.582900000000e-08, + 4.618120000000e-08, + 4.653550000000e-08, + 4.689190000000e-08,  \
+ 4.725040000000e-08, + 4.761100000000e-08, + 4.797380000000e-08, + 4.833880000000e-08, + 4.870590000000e-08 ]

.param id_pred_data_vg0.13=[ \
+ 7.961099299791e-09, + 1.349756416857e-08, + 1.735140926939e-08, + 2.004281441259e-08, + 2.193568917619e-08,  \
+ 2.328397613383e-08, + 2.426447622383e-08, + 2.499994707250e-08, + 2.557515159651e-08, + 2.604829489883e-08,  \
+ 2.645884705998e-08, + 2.683318143681e-08, + 2.718873361118e-08, + 2.753620350404e-08, + 2.788211688198e-08,  \
+ 2.822974238370e-08, + 2.858047665200e-08, + 2.893406218618e-08, + 2.928972065774e-08, + 2.964603140754e-08,  \
+ 3.000138846687e-08, + 3.035410145458e-08, + 3.070279916528e-08, + 3.104602569692e-08, + 3.138285009641e-08,  \
+ 3.171243747602e-08, + 3.203426643950e-08, + 3.234808559682e-08, + 3.265403670127e-08, + 3.295220736277e-08,  \
+ 3.324318576858e-08, + 3.352753310537e-08, + 3.380591444113e-08, + 3.407934642041e-08, + 3.434832578364e-08,  \
+ 3.461413683681e-08, + 3.487743128971e-08, + 3.513930323606e-08, + 3.540049448247e-08, + 3.566180453163e-08,  \
+ 3.592396190299e-08, + 3.618770136882e-08, + 3.645356294157e-08, + 3.672217872008e-08, + 3.699397908008e-08,  \
+ 3.726921534053e-08, + 3.754823005409e-08, + 3.783132569879e-08, + 3.811876347015e-08, + 3.841040907560e-08,  \
+ 3.870637144132e-08, + 3.900679985236e-08, + 3.931143872649e-08, + 3.962029680338e-08, + 3.993319026563e-08,  \
+ 4.024983695672e-08, + 4.057021683934e-08, + 4.089397307894e-08, + 4.122071210588e-08, + 4.155033224151e-08,  \
+ 4.188245718240e-08, + 4.221675780514e-08, + 4.255288153843e-08, + 4.289044682082e-08, + 4.322911983934e-08,  \
+ 4.356854802268e-08, + 4.390834860146e-08, + 4.424820218674e-08, + 4.458767499216e-08, + 4.492639789078e-08,  \
+ 4.526389297155e-08, + 4.560000888887e-08, + 4.593431398803e-08, + 4.626635757177e-08, + 4.659584718070e-08,  \
+ 4.692238093185e-08, + 4.724581970095e-08, + 4.756555256336e-08, + 4.788158470603e-08, + 4.819327728001e-08 ]

* Data table for Id-Vd at Vg = 0.14V
.param vd_data_vg0.14=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.14=[ \
+ 1.168790000000e-08, + 1.975940000000e-08, + 2.529830000000e-08, + 2.909780000000e-08, + 3.176760000000e-08,  \
+ 3.372640000000e-08, + 3.521550000000e-08, + 3.637710000000e-08, + 3.731070000000e-08, + 3.808810000000e-08,  \
+ 3.875900000000e-08, + 3.935690000000e-08, + 3.990390000000e-08, + 4.041480000000e-08, + 4.089960000000e-08,  \
+ 4.136520000000e-08, + 4.181630000000e-08, + 4.225660000000e-08, + 4.268860000000e-08, + 4.311420000000e-08,  \
+ 4.353490000000e-08, + 4.395180000000e-08, + 4.436590000000e-08, + 4.477780000000e-08, + 4.518810000000e-08,  \
+ 4.559740000000e-08, + 4.600610000000e-08, + 4.641440000000e-08, + 4.682260000000e-08, + 4.723110000000e-08,  \
+ 4.764000000000e-08, + 4.804960000000e-08, + 4.845990000000e-08, + 4.887120000000e-08, + 4.928350000000e-08,  \
+ 4.969700000000e-08, + 5.011180000000e-08, + 5.052790000000e-08, + 5.094560000000e-08, + 5.136480000000e-08,  \
+ 5.178560000000e-08, + 5.220810000000e-08, + 5.263240000000e-08, + 5.305850000000e-08, + 5.348650000000e-08,  \
+ 5.391640000000e-08, + 5.434830000000e-08, + 5.478230000000e-08, + 5.521830000000e-08, + 5.565640000000e-08,  \
+ 5.609670000000e-08, + 5.653920000000e-08, + 5.698390000000e-08, + 5.743090000000e-08, + 5.788020000000e-08,  \
+ 5.833190000000e-08, + 5.878590000000e-08, + 5.924230000000e-08, + 5.970120000000e-08, + 6.016250000000e-08,  \
+ 6.062630000000e-08, + 6.109270000000e-08, + 6.156150000000e-08, + 6.203300000000e-08, + 6.250710000000e-08,  \
+ 6.298380000000e-08, + 6.346310000000e-08, + 6.394520000000e-08, + 6.442990000000e-08, + 6.491730000000e-08,  \
+ 6.540760000000e-08, + 6.590060000000e-08, + 6.639630000000e-08, + 6.689500000000e-08, + 6.739640000000e-08,  \
+ 6.790070000000e-08, + 6.840800000000e-08, + 6.891810000000e-08, + 6.943120000000e-08, + 6.994720000000e-08 ]

.param id_pred_data_vg0.14=[ \
+ 1.146998670265e-08, + 1.949491434061e-08, + 2.510861577321e-08, + 2.904286247940e-08, + 3.181422414400e-08,  \
+ 3.378641622476e-08, + 3.521495955283e-08, + 3.627864316513e-08, + 3.710213064778e-08, + 3.777169581554e-08,  \
+ 3.834654052071e-08, + 3.886673766829e-08, + 3.935887576745e-08, + 3.983976114341e-08, + 4.031965374907e-08,  \
+ 4.080428880116e-08, + 4.129592809932e-08, + 4.179474558441e-08, + 4.229965540503e-08, + 4.280855421257e-08,  \
+ 4.331908186828e-08, + 4.382857440532e-08, + 4.433464269482e-08, + 4.483500674723e-08, + 4.532769892762e-08,  \
+ 4.581129530834e-08, + 4.628450071209e-08, + 4.674660942783e-08, + 4.719734292280e-08, + 4.763680436781e-08,  \
+ 4.806501635812e-08, + 4.848289336223e-08, + 4.889109234796e-08, + 4.929081541150e-08, + 4.968307578679e-08,  \
+ 5.006908168070e-08, + 5.045022945183e-08, + 5.082767017939e-08, + 5.120273740999e-08, + 5.157660893929e-08,  \
+ 5.195045574169e-08, + 5.232536580024e-08, + 5.270225258869e-08, + 5.308199206411e-08, + 5.346539531104e-08,  \
+ 5.385310942074e-08, + 5.424562367295e-08, + 5.464340233630e-08, + 5.504681780621e-08, + 5.545602732582e-08,  \
+ 5.587149708219e-08, + 5.629280764197e-08, + 5.672044181892e-08, + 5.715408050833e-08, + 5.759358181479e-08,  \
+ 5.803875296806e-08, + 5.848945498599e-08, + 5.894530133332e-08, + 5.940585197095e-08, + 5.987083682157e-08,  \
+ 6.033996321264e-08, + 6.081265794933e-08, + 6.128842393593e-08, + 6.176683655212e-08, + 6.224744133476e-08,  \
+ 6.272949562458e-08, + 6.321295266787e-08, + 6.369687298502e-08, + 6.418077909132e-08, + 6.466415385376e-08,  \
+ 6.514669451008e-08, + 6.562757505435e-08, + 6.610643502825e-08, + 6.658239641411e-08, + 6.705541721885e-08,  \
+ 6.752481283456e-08, + 6.799013434033e-08, + 6.845037816561e-08, + 6.890583350128e-08, + 6.935531473573e-08 ]

* Data table for Id-Vd at Vg = 0.15V
.param vd_data_vg0.15=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.15=[ \
+ 1.686830000000e-08, + 2.855550000000e-08, + 3.659350000000e-08, + 4.211440000000e-08, + 4.599460000000e-08,  \
+ 4.884020000000e-08, + 5.100170000000e-08, + 5.268640000000e-08, + 5.403840000000e-08, + 5.516210000000e-08,  \
+ 5.613010000000e-08, + 5.699100000000e-08, + 5.777730000000e-08, + 5.851040000000e-08, + 5.920510000000e-08,  \
+ 5.987130000000e-08, + 6.051620000000e-08, + 6.114490000000e-08, + 6.176120000000e-08, + 6.236790000000e-08,  \
+ 6.296720000000e-08, + 6.356070000000e-08, + 6.414970000000e-08, + 6.473530000000e-08, + 6.531850000000e-08,  \
+ 6.589980000000e-08, + 6.647990000000e-08, + 6.705930000000e-08, + 6.763840000000e-08, + 6.821750000000e-08,  \
+ 6.879700000000e-08, + 6.937720000000e-08, + 6.995830000000e-08, + 7.054050000000e-08, + 7.112400000000e-08,  \
+ 7.170900000000e-08, + 7.229560000000e-08, + 7.288400000000e-08, + 7.347420000000e-08, + 7.406650000000e-08,  \
+ 7.466090000000e-08, + 7.525750000000e-08, + 7.585650000000e-08, + 7.645780000000e-08, + 7.706170000000e-08,  \
+ 7.766800000000e-08, + 7.827710000000e-08, + 7.888880000000e-08, + 7.950320000000e-08, + 8.012050000000e-08,  \
+ 8.074070000000e-08, + 8.136380000000e-08, + 8.198990000000e-08, + 8.261900000000e-08, + 8.325120000000e-08,  \
+ 8.388660000000e-08, + 8.452510000000e-08, + 8.516680000000e-08, + 8.581180000000e-08, + 8.646010000000e-08,  \
+ 8.711180000000e-08, + 8.776680000000e-08, + 8.842520000000e-08, + 8.908720000000e-08, + 8.975260000000e-08,  \
+ 9.042150000000e-08, + 9.109400000000e-08, + 9.177010000000e-08, + 9.244980000000e-08, + 9.313320000000e-08,  \
+ 9.382020000000e-08, + 9.451100000000e-08, + 9.520560000000e-08, + 9.590400000000e-08, + 9.660610000000e-08,  \
+ 9.731220000000e-08, + 9.802210000000e-08, + 9.873590000000e-08, + 9.945360000000e-08, + 1.001750000000e-07 ]

.param id_pred_data_vg0.15=[ \
+ 1.648744500926e-08, + 2.810066689563e-08, + 3.627082378443e-08, + 4.202117906971e-08, + 4.608139363427e-08,  \
+ 4.896995619674e-08, + 5.105474315314e-08, + 5.259542376734e-08, + 5.377482011681e-08, + 5.472063548950e-08,  \
+ 5.552159393574e-08, + 5.623829679280e-08, + 5.691141325315e-08, + 5.756754319464e-08, + 5.822304132153e-08,  \
+ 5.888731266168e-08, + 5.956484017133e-08, + 6.025651146047e-08, + 6.096107455278e-08, + 6.167583705974e-08,  \
+ 6.239714792855e-08, + 6.312145558240e-08, + 6.384462892584e-08, + 6.456315077230e-08, + 6.527381657406e-08,  \
+ 6.597379979212e-08, + 6.666099352515e-08, + 6.733354211974e-08, + 6.799061921470e-08, + 6.863174775162e-08,  \
+ 6.925700247962e-08, + 6.986665539443e-08, + 7.046167382896e-08, + 7.104344888376e-08, + 7.161284472090e-08,  \
+ 7.217198742637e-08, + 7.272249746393e-08, + 7.326600950819e-08, + 7.380447485161e-08, + 7.433940822921e-08,  \
+ 7.487281877161e-08, + 7.540618327084e-08, + 7.594098065056e-08, + 7.647875463590e-08, + 7.702042523761e-08,  \
+ 7.756726802199e-08, + 7.812010281327e-08, + 7.868012289691e-08, + 7.924738667953e-08, + 7.982271910123e-08,  \
+ 8.040632309303e-08, + 8.099850617782e-08, + 8.159950155573e-08, + 8.220915788115e-08, + 8.282734356158e-08,  \
+ 8.345402306986e-08, + 8.408878031219e-08, + 8.473136887233e-08, + 8.538125626956e-08, + 8.603798846707e-08,  \
+ 8.670122781496e-08, + 8.736993805769e-08, + 8.804406675722e-08, + 8.872236321622e-08, + 8.940469413687e-08,  \
+ 9.008984449110e-08, + 9.077732741503e-08, + 9.146642526048e-08, + 9.215628750781e-08, + 9.284618727179e-08,  \
+ 9.353537620882e-08, + 9.422275184079e-08, + 9.490809432577e-08, + 9.559005178517e-08, + 9.626804953200e-08,  \
+ 9.694138782379e-08, + 9.760932513814e-08, + 9.827072489088e-08, + 9.892544866830e-08, + 9.957217343981e-08 ]

* Data table for Id-Vd at Vg = 0.16V
.param vd_data_vg0.16=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.16=[ \
+ 2.423110000000e-08, + 4.109760000000e-08, + 5.273540000000e-08, + 6.074440000000e-08, + 6.637600000000e-08,  \
+ 7.050410000000e-08, + 7.363770000000e-08, + 7.607750000000e-08, + 7.803240000000e-08, + 7.965400000000e-08,  \
+ 8.104760000000e-08, + 8.228430000000e-08, + 8.341130000000e-08, + 8.446020000000e-08, + 8.545220000000e-08,  \
+ 8.640230000000e-08, + 8.732070000000e-08, + 8.821510000000e-08, + 8.909080000000e-08, + 8.995210000000e-08,  \
+ 9.080210000000e-08, + 9.164320000000e-08, + 9.247740000000e-08, + 9.330630000000e-08, + 9.413120000000e-08,  \
+ 9.495300000000e-08, + 9.577260000000e-08, + 9.659080000000e-08, + 9.740810000000e-08, + 9.822520000000e-08,  \
+ 9.904250000000e-08, + 9.986030000000e-08, + 1.006790000000e-07, + 1.014990000000e-07, + 1.023210000000e-07,  \
+ 1.031440000000e-07, + 1.039690000000e-07, + 1.047960000000e-07, + 1.056260000000e-07, + 1.064590000000e-07,  \
+ 1.072940000000e-07, + 1.081320000000e-07, + 1.089720000000e-07, + 1.098160000000e-07, + 1.106640000000e-07,  \
+ 1.115140000000e-07, + 1.123680000000e-07, + 1.132250000000e-07, + 1.140870000000e-07, + 1.149510000000e-07,  \
+ 1.158200000000e-07, + 1.166920000000e-07, + 1.175680000000e-07, + 1.184490000000e-07, + 1.193330000000e-07,  \
+ 1.202220000000e-07, + 1.211140000000e-07, + 1.220110000000e-07, + 1.229120000000e-07, + 1.238180000000e-07,  \
+ 1.247280000000e-07, + 1.256420000000e-07, + 1.265610000000e-07, + 1.274850000000e-07, + 1.284130000000e-07,  \
+ 1.293460000000e-07, + 1.302840000000e-07, + 1.312260000000e-07, + 1.321730000000e-07, + 1.331250000000e-07,  \
+ 1.340820000000e-07, + 1.350440000000e-07, + 1.360110000000e-07, + 1.369820000000e-07, + 1.379590000000e-07,  \
+ 1.389410000000e-07, + 1.399280000000e-07, + 1.409210000000e-07, + 1.419180000000e-07, + 1.429210000000e-07 ]

.param id_pred_data_vg0.16=[ \
+ 2.361348151680e-08, + 4.037383405375e-08, + 5.224448159424e-08, + 6.064481567591e-08, + 6.659748237325e-08,  \
+ 7.083703394528e-08, + 7.388982112388e-08, + 7.613099114678e-08, + 7.782760803821e-08, + 7.916808044683e-08,  \
+ 8.028475690480e-08, + 8.126902457661e-08, + 8.218355389999e-08, + 8.306962399729e-08, + 8.395375061809e-08,  \
+ 8.485144462611e-08, + 8.577091534789e-08, + 8.671494242662e-08, + 8.768253906055e-08, + 8.867025940162e-08,  \
+ 8.967357587153e-08, + 9.068683141322e-08, + 9.170447015094e-08, + 9.272079296352e-08, + 9.373076181873e-08,  \
+ 9.472968486079e-08, + 9.571384197216e-08, + 9.668025427345e-08, + 9.762658891077e-08, + 9.855168627837e-08,  \
+ 9.945464711336e-08, + 1.003355737339e-07, + 1.011953938246e-07, + 1.020351976422e-07, + 1.028563261229e-07,  \
+ 1.036613866745e-07, + 1.044521857807e-07, + 1.052311301919e-07, + 1.060009876142e-07, + 1.067638891072e-07,  \
+ 1.075224699321e-07, + 1.082792215357e-07, + 1.090363559797e-07, + 1.097954964280e-07, + 1.105594336082e-07,  \
+ 1.113291119736e-07, + 1.121063178289e-07, + 1.128924282057e-07, + 1.136884698383e-07, + 1.144951653487e-07,  \
+ 1.153133550247e-07, + 1.161434630603e-07, + 1.169860270522e-07, + 1.178408462010e-07, + 1.187080705733e-07,  \
+ 1.195874085624e-07, + 1.204787254494e-07, + 1.213816929635e-07, + 1.222956503000e-07, + 1.232199792867e-07,  \
+ 1.241538677732e-07, + 1.250965320310e-07, + 1.260474425635e-07, + 1.270053235203e-07, + 1.279693734091e-07,  \
+ 1.289386329972e-07, + 1.299116622988e-07, + 1.308878410100e-07, + 1.318657264449e-07, + 1.328444156456e-07,  \
+ 1.338227180270e-07, + 1.347994714251e-07, + 1.357734808494e-07, + 1.367433355881e-07, + 1.377082341492e-07,  \
+ 1.386666616554e-07, + 1.396178367941e-07, + 1.405601378224e-07, + 1.414930855503e-07, + 1.424147171747e-07 ]

* Data table for Id-Vd at Vg = 0.17V
.param vd_data_vg0.17=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.17=[ \
+ 3.458240000000e-08, + 5.881010000000e-08, + 7.560430000000e-08, + 8.719530000000e-08, + 9.535320000000e-08,  \
+ 1.013310000000e-07, + 1.058650000000e-07, + 1.093920000000e-07, + 1.122130000000e-07, + 1.145470000000e-07,  \
+ 1.165480000000e-07, + 1.183180000000e-07, + 1.199280000000e-07, + 1.214220000000e-07, + 1.228330000000e-07,  \
+ 1.241810000000e-07, + 1.254820000000e-07, + 1.267480000000e-07, + 1.279860000000e-07, + 1.292020000000e-07,  \
+ 1.304000000000e-07, + 1.315850000000e-07, + 1.327600000000e-07, + 1.339260000000e-07, + 1.350850000000e-07,  \
+ 1.362400000000e-07, + 1.373900000000e-07, + 1.385380000000e-07, + 1.396850000000e-07, + 1.408300000000e-07,  \
+ 1.419740000000e-07, + 1.431190000000e-07, + 1.442650000000e-07, + 1.454120000000e-07, + 1.465610000000e-07,  \
+ 1.477110000000e-07, + 1.488640000000e-07, + 1.500190000000e-07, + 1.511780000000e-07, + 1.523390000000e-07,  \
+ 1.535040000000e-07, + 1.546720000000e-07, + 1.558440000000e-07, + 1.570190000000e-07, + 1.581990000000e-07,  \
+ 1.593830000000e-07, + 1.605720000000e-07, + 1.617640000000e-07, + 1.629620000000e-07, + 1.641640000000e-07,  \
+ 1.653710000000e-07, + 1.665830000000e-07, + 1.678000000000e-07, + 1.690220000000e-07, + 1.702500000000e-07,  \
+ 1.714820000000e-07, + 1.727200000000e-07, + 1.739640000000e-07, + 1.752130000000e-07, + 1.764680000000e-07,  \
+ 1.777290000000e-07, + 1.789950000000e-07, + 1.802670000000e-07, + 1.815450000000e-07, + 1.828290000000e-07,  \
+ 1.841200000000e-07, + 1.854160000000e-07, + 1.867190000000e-07, + 1.880270000000e-07, + 1.893420000000e-07,  \
+ 1.906640000000e-07, + 1.919920000000e-07, + 1.933260000000e-07, + 1.946670000000e-07, + 1.960140000000e-07,  \
+ 1.973680000000e-07, + 1.987290000000e-07, + 2.000960000000e-07, + 2.014700000000e-07, + 2.028520000000e-07 ]

.param id_pred_data_vg0.17=[ \
+ 3.362896677572e-08, + 5.770816642325e-08, + 7.489924200854e-08, + 8.714865543880e-08, + 9.587531621946e-08,  \
+ 1.021099569698e-07, + 1.065985827609e-07, + 1.098793109122e-07, + 1.123392758018e-07, + 1.142550900113e-07,  \
+ 1.158222596587e-07, + 1.171790472654e-07, + 1.184208628047e-07, + 1.196119274027e-07, + 1.207944080761e-07,  \
+ 1.219947716891e-07, + 1.232270409446e-07, + 1.244976908765e-07, + 1.258070636823e-07, + 1.271517135137e-07,  \
+ 1.285259702399e-07, + 1.299219695738e-07, + 1.313317750373e-07, + 1.327476411461e-07, + 1.341612403394e-07,  \
+ 1.355658207558e-07, + 1.369552995811e-07, + 1.383243943565e-07, + 1.396688992372e-07, + 1.409861965840e-07,  \
+ 1.422741601687e-07, + 1.435325793864e-07, + 1.447614704375e-07, + 1.459612951749e-07, + 1.471347971460e-07,  \
+ 1.482831726207e-07, + 1.494099598176e-07, + 1.505180023287e-07, + 1.516109298905e-07, + 1.526915980321e-07,  \
+ 1.537640471838e-07, + 1.548310450517e-07, + 1.558962787840e-07, + 1.569626749642e-07, + 1.580335350582e-07,  \
+ 1.591109497667e-07, + 1.601971459309e-07, + 1.612943106011e-07, + 1.624042312187e-07, + 1.635288384705e-07,  \
+ 1.646686831691e-07, + 1.658246708303e-07, + 1.669977029906e-07, + 1.681879621174e-07, + 1.693959731597e-07,  \
+ 1.706208399810e-07, + 1.718630323921e-07, + 1.731217071210e-07, + 1.743961456668e-07, + 1.756859489888e-07,  \
+ 1.769899645865e-07, + 1.783067415317e-07, + 1.796359285322e-07, + 1.809756759030e-07, + 1.823239955456e-07,  \
+ 1.836809497036e-07, + 1.850438013662e-07, + 1.864114938144e-07, + 1.877825221186e-07, + 1.891545764465e-07,  \
+ 1.905268402425e-07, + 1.918969815051e-07, + 1.932636510560e-07, + 1.946248613649e-07, + 1.959793181072e-07,  \
+ 1.973241023734e-07, + 1.986588620184e-07, + 1.999811371434e-07, + 2.012895075154e-07, + 2.025816684181e-07 ]

* Data table for Id-Vd at Vg = 0.18V
.param vd_data_vg0.18=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.18=[ \
+ 4.892220000000e-08, + 8.349890000000e-08, + 1.076220000000e-07, + 1.243410000000e-07, + 1.361270000000e-07,  \
+ 1.447610000000e-07, + 1.513050000000e-07, + 1.563890000000e-07, + 1.604480000000e-07, + 1.637980000000e-07,  \
+ 1.666590000000e-07, + 1.691840000000e-07, + 1.714710000000e-07, + 1.735890000000e-07, + 1.755820000000e-07,  \
+ 1.774840000000e-07, + 1.793160000000e-07, + 1.810940000000e-07, + 1.828310000000e-07, + 1.845350000000e-07,  \
+ 1.862120000000e-07, + 1.878690000000e-07, + 1.895100000000e-07, + 1.911370000000e-07, + 1.927530000000e-07,  \
+ 1.943620000000e-07, + 1.959630000000e-07, + 1.975600000000e-07, + 1.991540000000e-07, + 2.007450000000e-07,  \
+ 2.023340000000e-07, + 2.039230000000e-07, + 2.055120000000e-07, + 2.071020000000e-07, + 2.086930000000e-07,  \
+ 2.102860000000e-07, + 2.118820000000e-07, + 2.134800000000e-07, + 2.150820000000e-07, + 2.166870000000e-07,  \
+ 2.182960000000e-07, + 2.199090000000e-07, + 2.215270000000e-07, + 2.231490000000e-07, + 2.247760000000e-07,  \
+ 2.264080000000e-07, + 2.280460000000e-07, + 2.296890000000e-07, + 2.313380000000e-07, + 2.329930000000e-07,  \
+ 2.346530000000e-07, + 2.363200000000e-07, + 2.379930000000e-07, + 2.396730000000e-07, + 2.413590000000e-07,  \
+ 2.430520000000e-07, + 2.447510000000e-07, + 2.464580000000e-07, + 2.481720000000e-07, + 2.498920000000e-07,  \
+ 2.516200000000e-07, + 2.533560000000e-07, + 2.550980000000e-07, + 2.568480000000e-07, + 2.586060000000e-07,  \
+ 2.603720000000e-07, + 2.621450000000e-07, + 2.639260000000e-07, + 2.657150000000e-07, + 2.675120000000e-07,  \
+ 2.693170000000e-07, + 2.711300000000e-07, + 2.729520000000e-07, + 2.747820000000e-07, + 2.766200000000e-07,  \
+ 2.784660000000e-07, + 2.803210000000e-07, + 2.821840000000e-07, + 2.840560000000e-07, + 2.859370000000e-07 ]

.param id_pred_data_vg0.18=[ \
+ 4.749799700221e-08, + 8.184872058337e-08, + 1.066047593667e-07, + 1.243966380571e-07, + 1.371651592308e-07,  \
+ 1.463373337174e-07, + 1.529590781502e-07, + 1.577928196639e-07, + 1.613942515633e-07, + 1.641640210437e-07,  \
+ 1.663911734795e-07, + 1.682807851466e-07, + 1.699775623365e-07, + 1.715809662528e-07, + 1.731582642606e-07,  \
+ 1.747517853801e-07, + 1.763870307059e-07, + 1.780772367965e-07, + 1.798253975949e-07, + 1.816297526602e-07,  \
+ 1.834830646885e-07, + 1.853765900250e-07, + 1.872991833807e-07, + 1.892397176562e-07, + 1.911868565685e-07,  \
+ 1.931304416303e-07, + 1.950604286094e-07, + 1.969698155335e-07, + 1.988505937334e-07, + 2.006986960623e-07,  \
+ 2.025097461456e-07, + 2.042820597126e-07, + 2.060145590121e-07, + 2.077076146634e-07, + 2.093631621847e-07,  \
+ 2.109833485520e-07, + 2.125711858980e-07, + 2.141308891623e-07, + 2.156669876285e-07, + 2.171833330067e-07,  \
+ 2.186847467556e-07, + 2.201762015375e-07, + 2.216622647211e-07, + 2.231468215541e-07, + 2.246345189860e-07,  \
+ 2.261286613248e-07, + 2.276332975271e-07, + 2.291510008945e-07, + 2.306847528644e-07, + 2.322365588725e-07,  \
+ 2.338087116982e-07, + 2.354026810281e-07, + 2.370188590817e-07, + 2.386583372527e-07, + 2.403220719316e-07,  \
+ 2.420092459943e-07, + 2.437197929339e-07, + 2.454534734397e-07, + 2.472092134553e-07, + 2.489859923571e-07,  \
+ 2.507828870080e-07, + 2.525978470658e-07, + 2.544296242490e-07, + 2.562760892033e-07, + 2.581359652254e-07,  \
+ 2.600065425895e-07, + 2.618862416170e-07, + 2.637720785970e-07, + 2.656627029296e-07, + 2.675548017805e-07,  \
+ 2.694462267527e-07, + 2.713344633776e-07, + 2.732176199061e-07, + 2.750924062411e-07, + 2.769566549432e-07,  \
+ 2.788071037685e-07, + 2.806422043022e-07, + 2.824589688544e-07, + 2.842551333515e-07, + 2.860272616090e-07 ]

* Data table for Id-Vd at Vg = 0.19V
.param vd_data_vg0.19=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.19=[ \
+ 6.840530000000e-08, + 1.173190000000e-07, + 1.517480000000e-07, + 1.757520000000e-07, + 1.927150000000e-07,  \
+ 2.051410000000e-07, + 2.145540000000e-07, + 2.218590000000e-07, + 2.276780000000e-07, + 2.324640000000e-07,  \
+ 2.365380000000e-07, + 2.401160000000e-07, + 2.433460000000e-07, + 2.463260000000e-07, + 2.491240000000e-07,  \
+ 2.517840000000e-07, + 2.543410000000e-07, + 2.568180000000e-07, + 2.592330000000e-07, + 2.615980000000e-07,  \
+ 2.639230000000e-07, + 2.662170000000e-07, + 2.684840000000e-07, + 2.707310000000e-07, + 2.729620000000e-07,  \
+ 2.751780000000e-07, + 2.773840000000e-07, + 2.795820000000e-07, + 2.817720000000e-07, + 2.839580000000e-07,  \
+ 2.861400000000e-07, + 2.883200000000e-07, + 2.904990000000e-07, + 2.926780000000e-07, + 2.948570000000e-07,  \
+ 2.970370000000e-07, + 2.992200000000e-07, + 3.014050000000e-07, + 3.035930000000e-07, + 3.057850000000e-07,  \
+ 3.079810000000e-07, + 3.101820000000e-07, + 3.123880000000e-07, + 3.145990000000e-07, + 3.168150000000e-07,  \
+ 3.190380000000e-07, + 3.212660000000e-07, + 3.235020000000e-07, + 3.257430000000e-07, + 3.279920000000e-07,  \
+ 3.302480000000e-07, + 3.325120000000e-07, + 3.347830000000e-07, + 3.370620000000e-07, + 3.393490000000e-07,  \
+ 3.416430000000e-07, + 3.439470000000e-07, + 3.462580000000e-07, + 3.485780000000e-07, + 3.509070000000e-07,  \
+ 3.532450000000e-07, + 3.555910000000e-07, + 3.579470000000e-07, + 3.603120000000e-07, + 3.626860000000e-07,  \
+ 3.650700000000e-07, + 3.674630000000e-07, + 3.698660000000e-07, + 3.722780000000e-07, + 3.747010000000e-07,  \
+ 3.771330000000e-07, + 3.795750000000e-07, + 3.820280000000e-07, + 3.844910000000e-07, + 3.869640000000e-07,  \
+ 3.894470000000e-07, + 3.919410000000e-07, + 3.944450000000e-07, + 3.969600000000e-07, + 3.994860000000e-07 ]

.param id_pred_data_vg0.19=[ \
+ 6.633278644586e-08, + 1.148444607679e-07, + 1.501863380327e-07, + 1.758481448633e-07, + 1.944390760400e-07,  \
+ 2.079014166156e-07, + 2.176764655815e-07, + 2.248303098895e-07, + 2.301471704413e-07, + 2.342020252399e-07,  \
+ 2.374140058237e-07, + 2.400854555162e-07, + 2.424329375117e-07, + 2.446080361551e-07, + 2.467156889452e-07,  \
+ 2.488254176569e-07, + 2.509804676265e-07, + 2.532054872972e-07, + 2.555107926128e-07, + 2.578971816547e-07,  \
+ 2.603583311611e-07, + 2.628841889418e-07, + 2.654612262631e-07, + 2.680737270566e-07, + 2.707083410769e-07,  \
+ 2.733489782258e-07, + 2.759826952570e-07, + 2.785970218611e-07, + 2.811821605064e-07, + 2.837294005076e-07,  \
+ 2.862323503905e-07, + 2.886864422180e-07, + 2.910900866482e-07, + 2.934411520528e-07, + 2.957414210414e-07,  \
+ 2.979933765346e-07, + 3.001999806429e-07, + 3.023663145996e-07, + 3.044961744081e-07, + 3.065967121074e-07,  \
+ 3.086741804736e-07, + 3.107337329311e-07, + 3.127811902459e-07, + 3.148240489281e-07, + 3.168670190234e-07,  \
+ 3.189150561411e-07, + 3.209745989352e-07, + 3.230493530282e-07, + 3.251414761962e-07, + 3.272575099800e-07,  \
+ 3.293975208862e-07, + 3.315666367598e-07, + 3.337634581158e-07, + 3.359913716849e-07, + 3.382494242032e-07,  \
+ 3.405396500966e-07, + 3.428606083844e-07, + 3.452119403846e-07, + 3.475927178442e-07, + 3.500015168356e-07,  \
+ 3.524363251017e-07, + 3.548952497567e-07, + 3.573768276510e-07, + 3.598777402658e-07, + 3.623951101872e-07,  \
+ 3.649268808203e-07, + 3.674690623257e-07, + 3.700192155520e-07, + 3.725732716475e-07, + 3.751284282316e-07,  \
+ 3.776812565093e-07, + 3.802282571996e-07, + 3.827660492561e-07, + 3.852896372791e-07, + 3.877967600374e-07,  \
+ 3.902827870661e-07, + 3.927440809548e-07, + 3.951783958200e-07, + 3.975806293965e-07, + 3.999474756711e-07 ]

* Data table for Id-Vd at Vg = 0.20V
.param vd_data_vg0.20=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.20=[ \
+ 9.423290000000e-08, + 1.626270000000e-07, + 2.113360000000e-07, + 2.455780000000e-07, + 2.698700000000e-07,  \
+ 2.876720000000e-07, + 3.011490000000e-07, + 3.115980000000e-07, + 3.199010000000e-07, + 3.267040000000e-07,  \
+ 3.324680000000e-07, + 3.375060000000e-07, + 3.420330000000e-07, + 3.461910000000e-07, + 3.500790000000e-07,  \
+ 3.537650000000e-07, + 3.572970000000e-07, + 3.607100000000e-07, + 3.640290000000e-07, + 3.672730000000e-07,  \
+ 3.704580000000e-07, + 3.735940000000e-07, + 3.766900000000e-07, + 3.797540000000e-07, + 3.827910000000e-07,  \
+ 3.858070000000e-07, + 3.888040000000e-07, + 3.917870000000e-07, + 3.947590000000e-07, + 3.977210000000e-07,  \
+ 4.006750000000e-07, + 4.036250000000e-07, + 4.065700000000e-07, + 4.095130000000e-07, + 4.124550000000e-07,  \
+ 4.153970000000e-07, + 4.183390000000e-07, + 4.212830000000e-07, + 4.242300000000e-07, + 4.271790000000e-07,  \
+ 4.301330000000e-07, + 4.330910000000e-07, + 4.360540000000e-07, + 4.390220000000e-07, + 4.419960000000e-07,  \
+ 4.449770000000e-07, + 4.479650000000e-07, + 4.509590000000e-07, + 4.539610000000e-07, + 4.569710000000e-07,  \
+ 4.599890000000e-07, + 4.630160000000e-07, + 4.660510000000e-07, + 4.690950000000e-07, + 4.721480000000e-07,  \
+ 4.752100000000e-07, + 4.782830000000e-07, + 4.813650000000e-07, + 4.844560000000e-07, + 4.875590000000e-07,  \
+ 4.906710000000e-07, + 4.937940000000e-07, + 4.969280000000e-07, + 5.000720000000e-07, + 5.032280000000e-07,  \
+ 5.063940000000e-07, + 5.095720000000e-07, + 5.127620000000e-07, + 5.159620000000e-07, + 5.191750000000e-07,  \
+ 5.223990000000e-07, + 5.256360000000e-07, + 5.288840000000e-07, + 5.321440000000e-07, + 5.354170000000e-07,  \
+ 5.387020000000e-07, + 5.419990000000e-07, + 5.453090000000e-07, + 5.486320000000e-07, + 5.519670000000e-07 ]

.param id_pred_data_vg0.20=[ \
+ 9.130706530414e-08, + 1.589088060427e-07, + 2.087576285703e-07, + 2.453843990224e-07, + 2.722191993598e-07,  \
+ 2.918547852460e-07, + 3.062376254093e-07, + 3.168278999510e-07, + 3.247158906561e-07, + 3.307080305603e-07,  \
+ 3.354043860782e-07, + 3.392421967874e-07, + 3.425409090596e-07, + 3.455284740994e-07, + 3.483657906145e-07,  \
+ 3.511621980579e-07, + 3.539911836015e-07, + 3.568958300093e-07, + 3.599000649501e-07, + 3.630113724284e-07,  \
+ 3.662275798888e-07, + 3.695372902257e-07, + 3.729268053121e-07, + 3.763775475818e-07, + 3.798699879098e-07,  \
+ 3.833864002445e-07, + 3.869061231399e-07, + 3.904129289367e-07, + 3.938932138681e-07, + 3.973330422014e-07,  \
+ 4.007227460079e-07, + 4.040547719342e-07, + 4.073237789726e-07, + 4.105279163014e-07, + 4.136662994370e-07,  \
+ 4.167399174548e-07, + 4.197533257866e-07, + 4.227106660437e-07, + 4.256183808593e-07, + 4.284829628887e-07,  \
+ 4.313118495247e-07, + 4.341130625107e-07, + 4.368943473310e-07, + 4.396639496917e-07, + 4.424284043125e-07,  \
+ 4.451971085473e-07, + 4.479747792629e-07, + 4.507685480348e-07, + 4.535831226349e-07, + 4.564240612126e-07,  \
+ 4.592957157001e-07, + 4.621994116860e-07, + 4.651397352973e-07, + 4.681169116338e-07, + 4.711348594810e-07,  \
+ 4.741909333461e-07, + 4.772857744229e-07, + 4.804192190022e-07, + 4.835890632648e-07, + 4.867945108344e-07,  \
+ 4.900332481839e-07, + 4.933015611641e-07, + 4.965960442860e-07, + 4.999148222851e-07, + 5.032528548554e-07,  \
+ 5.066072958471e-07, + 5.099725410673e-07, + 5.133446688887e-07, + 5.167204818690e-07, + 5.200925500048e-07,  \
+ 5.234571796109e-07, + 5.268098584565e-07, + 5.301454820028e-07, + 5.334570437299e-07, + 5.367424478209e-07,  \
+ 5.399958467933e-07, + 5.432101278302e-07, + 5.463805416639e-07, + 5.495053812865e-07, + 5.525742380996e-07 ]

* Data table for Id-Vd at Vg = 0.21V
.param vd_data_vg0.21=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.21=[ \
+ 1.274660000000e-07, + 2.216860000000e-07, + 2.898030000000e-07, + 3.382250000000e-07, + 3.727770000000e-07,  \
+ 3.981260000000e-07, + 4.173120000000e-07, + 4.321700000000e-07, + 4.439490000000e-07, + 4.535590000000e-07,  \
+ 4.616560000000e-07, + 4.686930000000e-07, + 4.749800000000e-07, + 4.807240000000e-07, + 4.860710000000e-07,  \
+ 4.911180000000e-07, + 4.959370000000e-07, + 5.005790000000e-07, + 5.050810000000e-07, + 5.094710000000e-07,  \
+ 5.137700000000e-07, + 5.179960000000e-07, + 5.221620000000e-07, + 5.262770000000e-07, + 5.303500000000e-07,  \
+ 5.343890000000e-07, + 5.383990000000e-07, + 5.423850000000e-07, + 5.463510000000e-07, + 5.503000000000e-07,  \
+ 5.542360000000e-07, + 5.581610000000e-07, + 5.620780000000e-07, + 5.659880000000e-07, + 5.698930000000e-07,  \
+ 5.737950000000e-07, + 5.776950000000e-07, + 5.815940000000e-07, + 5.854940000000e-07, + 5.893960000000e-07,  \
+ 5.933000000000e-07, + 5.972070000000e-07, + 6.011180000000e-07, + 6.050340000000e-07, + 6.089560000000e-07,  \
+ 6.128840000000e-07, + 6.168180000000e-07, + 6.207590000000e-07, + 6.247080000000e-07, + 6.286650000000e-07,  \
+ 6.326300000000e-07, + 6.366050000000e-07, + 6.405880000000e-07, + 6.445810000000e-07, + 6.485840000000e-07,  \
+ 6.525980000000e-07, + 6.566210000000e-07, + 6.606560000000e-07, + 6.647010000000e-07, + 6.687580000000e-07,  \
+ 6.728270000000e-07, + 6.769070000000e-07, + 6.809990000000e-07, + 6.851030000000e-07, + 6.892200000000e-07,  \
+ 6.933490000000e-07, + 6.974910000000e-07, + 7.016460000000e-07, + 7.058140000000e-07, + 7.099950000000e-07,  \
+ 7.141890000000e-07, + 7.183980000000e-07, + 7.226190000000e-07, + 7.268550000000e-07, + 7.311050000000e-07,  \
+ 7.353680000000e-07, + 7.396460000000e-07, + 7.439380000000e-07, + 7.482450000000e-07, + 7.525670000000e-07 ]

.param id_pred_data_vg0.21=[ \
+ 1.235211311723e-07, + 2.161866723327e-07, + 2.854238300642e-07, + 3.369668775122e-07, + 3.752195880224e-07,  \
+ 4.035554866277e-07, + 4.245464970154e-07, + 4.401463957038e-07, + 4.518352898231e-07, + 4.607256414602e-07,  \
+ 4.676530761571e-07, + 4.732409979624e-07, + 4.779484288520e-07, + 4.821105585506e-07, + 4.859697924076e-07,  \
+ 4.896970131085e-07, + 4.934076446261e-07, + 4.971783573637e-07, + 5.010527388549e-07, + 5.050542768004e-07,  \
+ 5.091874118079e-07, + 5.134457569511e-07, + 5.178163564779e-07, + 5.222784602665e-07, + 5.268101403999e-07,  \
+ 5.313856081557e-07, + 5.359849114939e-07, + 5.405830506788e-07, + 5.451611991703e-07, + 5.497002234733e-07,  \
+ 5.541868415548e-07, + 5.586089537246e-07, + 5.629576889987e-07, + 5.672286101799e-07, + 5.714188546335e-07,  \
+ 5.755284837505e-07, + 5.795607603432e-07, + 5.835192973791e-07, + 5.874116459381e-07, + 5.912466804148e-07,  \
+ 5.950298861990e-07, + 5.987733334223e-07, + 6.024859578702e-07, + 6.061769272492e-07, + 6.098580968228e-07,  \
+ 6.135365015325e-07, + 6.172219877953e-07, + 6.209226012288e-07, + 6.246470763926e-07, + 6.283981974775e-07,  \
+ 6.321835974177e-07, + 6.360086672430e-07, + 6.398758625892e-07, + 6.437872571041e-07, + 6.477449574049e-07,  \
+ 6.517495785374e-07, + 6.558012637470e-07, + 6.598977142858e-07, + 6.640383128342e-07, + 6.682199455099e-07,  \
+ 6.724406330250e-07, + 6.766970454919e-07, + 6.809824742504e-07, + 6.852923252154e-07, + 6.896247498389e-07,  \
+ 6.939699801478e-07, + 6.983253274484e-07, + 7.026842058622e-07, + 7.070387232488e-07, + 7.113833930816e-07,  \
+ 7.157104494127e-07, + 7.200149775599e-07, + 7.242878666602e-07, + 7.285244828381e-07, + 7.327155628900e-07,  \
+ 7.368538535957e-07, + 7.409346437726e-07, + 7.449493182321e-07, + 7.488911086284e-07, + 7.527518846473e-07 ]

* Data table for Id-Vd at Vg = 0.22V
.param vd_data_vg0.22=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.22=[ \
+ 1.687960000000e-07, + 2.962440000000e-07, + 3.900970000000e-07, + 4.577830000000e-07, + 5.064870000000e-07,  \
+ 5.423090000000e-07, + 5.694210000000e-07, + 5.904030000000e-07, + 6.069940000000e-07, + 6.204690000000e-07,  \
+ 6.317530000000e-07, + 6.414950000000e-07, + 6.501380000000e-07, + 6.579870000000e-07, + 6.652510000000e-07,  \
+ 6.720740000000e-07, + 6.785600000000e-07, + 6.847830000000e-07, + 6.907990000000e-07, + 6.966480000000e-07,  \
+ 7.023610000000e-07, + 7.079640000000e-07, + 7.134750000000e-07, + 7.189090000000e-07, + 7.242790000000e-07,  \
+ 7.295950000000e-07, + 7.348650000000e-07, + 7.400970000000e-07, + 7.452960000000e-07, + 7.504670000000e-07,  \
+ 7.556150000000e-07, + 7.607440000000e-07, + 7.658560000000e-07, + 7.709540000000e-07, + 7.760420000000e-07,  \
+ 7.811210000000e-07, + 7.861930000000e-07, + 7.912600000000e-07, + 7.963240000000e-07, + 8.013860000000e-07,  \
+ 8.064470000000e-07, + 8.115090000000e-07, + 8.165730000000e-07, + 8.216400000000e-07, + 8.267100000000e-07,  \
+ 8.317840000000e-07, + 8.368640000000e-07, + 8.419500000000e-07, + 8.470420000000e-07, + 8.521420000000e-07,  \
+ 8.572500000000e-07, + 8.623660000000e-07, + 8.674910000000e-07, + 8.726250000000e-07, + 8.777690000000e-07,  \
+ 8.829230000000e-07, + 8.880880000000e-07, + 8.932640000000e-07, + 8.984510000000e-07, + 9.036500000000e-07,  \
+ 9.088610000000e-07, + 9.140850000000e-07, + 9.193200000000e-07, + 9.245690000000e-07, + 9.298310000000e-07,  \
+ 9.351060000000e-07, + 9.403950000000e-07, + 9.456980000000e-07, + 9.510150000000e-07, + 9.563460000000e-07,  \
+ 9.616920000000e-07, + 9.670520000000e-07, + 9.724270000000e-07, + 9.778170000000e-07, + 9.832220000000e-07,  \
+ 9.886430000000e-07, + 9.940790000000e-07, + 9.995310000000e-07, + 1.005000000000e-06, + 1.010500000000e-06 ]

.param id_pred_data_vg0.22=[ \
+ 1.638347202970e-07, + 2.884577588702e-07, + 3.828816807072e-07, + 4.541664384305e-07, + 5.078163667349e-07,  \
+ 5.481073276314e-07, + 5.783459801023e-07, + 6.010840661475e-07, + 6.182780316522e-07, + 6.314235179161e-07,  \
+ 6.416612313842e-07, + 6.498524453491e-07, + 6.566435104105e-07, + 6.625190872001e-07, + 6.678313411612e-07,  \
+ 6.728385051247e-07, + 6.777203680031e-07, + 6.826000935689e-07, + 6.875586632304e-07, + 6.926426522114e-07,  \
+ 6.978735677876e-07, + 7.032543271634e-07, + 7.087761514413e-07, + 7.144216397137e-07, + 7.201677476587e-07,  \
+ 7.259856283781e-07, + 7.318496068365e-07, + 7.377318434010e-07, + 7.436058103849e-07, + 7.494489636883e-07,  \
+ 7.552417423540e-07, + 7.609676686116e-07, + 7.666131068618e-07, + 7.721720339759e-07, + 7.776359893796e-07,  \
+ 7.830046524759e-07, + 7.882799445724e-07, + 7.934643554108e-07, + 7.985644401742e-07, + 8.035887731239e-07,  \
+ 8.085486456366e-07, + 8.134537574733e-07, + 8.183133172679e-07, + 8.231420042648e-07, + 8.279512371701e-07,  \
+ 8.327512728101e-07, + 8.375538516248e-07, + 8.423698636761e-07, + 8.472068896026e-07, + 8.520742653673e-07,  \
+ 8.569782153245e-07, + 8.619258233011e-07, + 8.669186286170e-07, + 8.719633297005e-07, + 8.770594547514e-07,  \
+ 8.822082781990e-07, + 8.874107584234e-07, + 8.926644977691e-07, + 8.979683570942e-07, + 9.033164360517e-07,  \
+ 9.087073760838e-07, + 9.141332475338e-07, + 9.195907318826e-07, + 9.250727453036e-07, + 9.305714229413e-07,  \
+ 9.360784702039e-07, + 9.415895783604e-07, + 9.470937675360e-07, + 9.525821496936e-07, + 9.580491337147e-07,  \
+ 9.634785374146e-07, + 9.688703266875e-07, + 9.742065662977e-07, + 9.794854759093e-07, + 9.846901320998e-07,  \
+ 9.898182497636e-07, + 9.948558283668e-07, + 9.997942424889e-07, + 1.004627417842e-06, + 1.009341485769e-06 ]

* Data table for Id-Vd at Vg = 0.23V
.param vd_data_vg0.23=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.23=[ \
+ 2.183400000000e-07, + 3.871040000000e-07, + 5.140750000000e-07, + 6.072940000000e-07, + 6.751480000000e-07,  \
+ 7.252770000000e-07, + 7.632530000000e-07, + 7.926320000000e-07, + 8.158120000000e-07, + 8.345510000000e-07,  \
+ 8.501400000000e-07, + 8.634970000000e-07, + 8.752560000000e-07, + 8.858570000000e-07, + 8.956010000000e-07,  \
+ 9.047000000000e-07, + 9.133040000000e-07, + 9.215230000000e-07, + 9.294350000000e-07, + 9.371010000000e-07,  \
+ 9.445670000000e-07, + 9.518670000000e-07, + 9.590310000000e-07, + 9.660790000000e-07, + 9.730300000000e-07,  \
+ 9.798980000000e-07, + 9.866960000000e-07, + 9.934340000000e-07, + 1.000100000000e-06, + 1.006800000000e-06,  \
+ 1.013400000000e-06, + 1.019900000000e-06, + 1.026500000000e-06, + 1.033000000000e-06, + 1.039500000000e-06,  \
+ 1.046000000000e-06, + 1.052400000000e-06, + 1.058900000000e-06, + 1.065300000000e-06, + 1.071800000000e-06,  \
+ 1.078200000000e-06, + 1.084600000000e-06, + 1.091000000000e-06, + 1.097500000000e-06, + 1.103900000000e-06,  \
+ 1.110300000000e-06, + 1.116700000000e-06, + 1.123200000000e-06, + 1.129600000000e-06, + 1.136000000000e-06,  \
+ 1.142500000000e-06, + 1.148900000000e-06, + 1.155400000000e-06, + 1.161800000000e-06, + 1.168300000000e-06,  \
+ 1.174800000000e-06, + 1.181300000000e-06, + 1.187800000000e-06, + 1.194300000000e-06, + 1.200800000000e-06,  \
+ 1.207300000000e-06, + 1.213900000000e-06, + 1.220400000000e-06, + 1.227000000000e-06, + 1.233600000000e-06,  \
+ 1.240200000000e-06, + 1.246800000000e-06, + 1.253400000000e-06, + 1.260100000000e-06, + 1.266700000000e-06,  \
+ 1.273400000000e-06, + 1.280100000000e-06, + 1.286800000000e-06, + 1.293500000000e-06, + 1.300200000000e-06,  \
+ 1.307000000000e-06, + 1.313700000000e-06, + 1.320500000000e-06, + 1.327300000000e-06, + 1.334100000000e-06 ]

.param id_pred_data_vg0.23=[ \
+ 2.127103289240e-07, + 3.768338865484e-07, + 5.029957719671e-07, + 5.996409527143e-07, + 6.734534963471e-07,  \
+ 7.297013689822e-07, + 7.725201703579e-07, + 8.051475015236e-07, + 8.301041543746e-07, + 8.493442692270e-07,  \
+ 8.643805631436e-07, + 8.763780715526e-07, + 8.862206095728e-07, + 8.945803529059e-07, + 9.019683602673e-07,  \
+ 9.087518265005e-07, + 9.152091706710e-07, + 9.215299269272e-07, + 9.278471088692e-07, + 9.342479643237e-07,  \
+ 9.407794505023e-07, + 9.474672515353e-07, + 9.543148189550e-07, + 9.613098882255e-07, + 9.684310953162e-07,  \
+ 9.756570034369e-07, + 9.829525379246e-07, + 9.902900001180e-07, + 9.976371893572e-07, + 1.004968362395e-06,  \
+ 1.012259122035e-06, + 1.019484407152e-06, + 1.026632498906e-06, + 1.033684466165e-06, + 1.040636561811e-06,  \
+ 1.047481200658e-06, + 1.054219721937e-06, + 1.060851577677e-06, + 1.067383152531e-06, + 1.073826388165e-06,  \
+ 1.080186341369e-06, + 1.086475222110e-06, + 1.092710447210e-06, + 1.098901484511e-06, + 1.105062563056e-06,  \
+ 1.111205269808e-06, + 1.117348315347e-06, + 1.123498841480e-06, + 1.129666786710e-06, + 1.135864522439e-06,  \
+ 1.142102075846e-06, + 1.148382552856e-06, + 1.154714261702e-06, + 1.161099207820e-06, + 1.167539858216e-06,  \
+ 1.174040189653e-06, + 1.180595413643e-06, + 1.187205507449e-06, + 1.193866594349e-06, + 1.200573797178e-06,  \
+ 1.207321895436e-06, + 1.214104627252e-06, + 1.220914052737e-06, + 1.227742613992e-06, + 1.234578661524e-06,  \
+ 1.241413556272e-06, + 1.248237703066e-06, + 1.255037664123e-06, + 1.261803917032e-06, + 1.268522748887e-06,  \
+ 1.275187438523e-06, + 1.281778313569e-06, + 1.288288566457e-06, + 1.294704979955e-06, + 1.301012588328e-06,  \
+ 1.307203197030e-06, + 1.313259804192e-06, + 1.319178518315e-06, + 1.324938942844e-06, + 1.330529084953e-06 ]

* Data table for Id-Vd at Vg = 0.24V
.param vd_data_vg0.24=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.24=[ \
+ 2.755740000000e-07, + 4.938470000000e-07, + 6.619870000000e-07, + 7.880430000000e-07, + 8.811830000000e-07,  \
+ 9.504910000000e-07, + 1.003100000000e-06, + 1.043800000000e-06, + 1.075900000000e-06, + 1.101800000000e-06,  \
+ 1.123100000000e-06, + 1.141200000000e-06, + 1.157100000000e-06, + 1.171200000000e-06, + 1.184100000000e-06,  \
+ 1.196100000000e-06, + 1.207400000000e-06, + 1.218000000000e-06, + 1.228300000000e-06, + 1.238200000000e-06,  \
+ 1.247800000000e-06, + 1.257100000000e-06, + 1.266300000000e-06, + 1.275200000000e-06, + 1.284100000000e-06,  \
+ 1.292800000000e-06, + 1.301400000000e-06, + 1.309900000000e-06, + 1.318300000000e-06, + 1.326700000000e-06,  \
+ 1.335000000000e-06, + 1.343200000000e-06, + 1.351400000000e-06, + 1.359600000000e-06, + 1.367700000000e-06,  \
+ 1.375800000000e-06, + 1.383900000000e-06, + 1.392000000000e-06, + 1.400000000000e-06, + 1.408000000000e-06,  \
+ 1.416000000000e-06, + 1.424000000000e-06, + 1.432000000000e-06, + 1.439900000000e-06, + 1.447900000000e-06,  \
+ 1.455800000000e-06, + 1.463800000000e-06, + 1.471800000000e-06, + 1.479700000000e-06, + 1.487700000000e-06,  \
+ 1.495600000000e-06, + 1.503600000000e-06, + 1.511500000000e-06, + 1.519500000000e-06, + 1.527500000000e-06,  \
+ 1.535500000000e-06, + 1.543400000000e-06, + 1.551400000000e-06, + 1.559400000000e-06, + 1.567400000000e-06,  \
+ 1.575500000000e-06, + 1.583500000000e-06, + 1.591500000000e-06, + 1.599600000000e-06, + 1.607600000000e-06,  \
+ 1.615700000000e-06, + 1.623800000000e-06, + 1.631900000000e-06, + 1.640000000000e-06, + 1.648100000000e-06,  \
+ 1.656300000000e-06, + 1.664400000000e-06, + 1.672600000000e-06, + 1.680800000000e-06, + 1.689000000000e-06,  \
+ 1.697200000000e-06, + 1.705400000000e-06, + 1.713700000000e-06, + 1.722000000000e-06, + 1.730200000000e-06 ]

.param id_pred_data_vg0.24=[ \
+ 2.701012999751e-07, + 4.815354259335e-07, + 6.464607758971e-07, + 7.746887422400e-07, + 8.741022611503e-07,  \
+ 9.510032032267e-07, + 1.010416999634e-06, + 1.056331748259e-06, + 1.091902831831e-06, + 1.119615080825e-06,  \
+ 1.141416660175e-06, + 1.158834238595e-06, + 1.173047648990e-06, + 1.184967077279e-06, + 1.195294589706e-06,  \
+ 1.204558648169e-06, + 1.213151390402e-06, + 1.221366810569e-06, + 1.229409863299e-06, + 1.237423748535e-06,  \
+ 1.245505613952e-06, + 1.253707914657e-06, + 1.262058467546e-06, + 1.270562606805e-06, + 1.279212028749e-06,  \
+ 1.287981449423e-06, + 1.296850309700e-06, + 1.305782298004e-06, + 1.314747846664e-06, + 1.323718606727e-06,  \
+ 1.332663218818e-06, + 1.341553579550e-06, + 1.350373781861e-06, + 1.359103853247e-06, + 1.367729191770e-06,  \
+ 1.376246127620e-06, + 1.384645240705e-06, + 1.392931862938e-06, + 1.401107269885e-06, + 1.409179185430e-06,  \
+ 1.417159055563e-06, + 1.425054956599e-06, + 1.432883389043e-06, + 1.440659716536e-06, + 1.448394300496e-06,  \
+ 1.456107906961e-06, + 1.463808710014e-06, + 1.471515461162e-06, + 1.479238426327e-06, + 1.486989503974e-06,  \
+ 1.494774710409e-06, + 1.502607583461e-06, + 1.510488846179e-06, + 1.518426861367e-06, + 1.526423068299e-06,  \
+ 1.534475068183e-06, + 1.542586558116e-06, + 1.550753127049e-06, + 1.558966216635e-06, + 1.567222443555e-06,  \
+ 1.575515832428e-06, + 1.583835278325e-06, + 1.592171647644e-06, + 1.600513351150e-06, + 1.608847969692e-06,  \
+ 1.617162529328e-06, + 1.625446075195e-06, + 1.633679166844e-06, + 1.641852384182e-06, + 1.649945102145e-06,  \
+ 1.657947893818e-06, + 1.665840063652e-06, + 1.673609879163e-06, + 1.681238159108e-06, + 1.688710312919e-06,  \
+ 1.696012959655e-06, + 1.703123593870e-06, + 1.710037740850e-06, + 1.716735191621e-06, + 1.723200875858e-06 ]

* Data table for Id-Vd at Vg = 0.25V
.param vd_data_vg0.25=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.25=[ \
+ 3.394150000000e-07, + 6.148470000000e-07, + 8.322910000000e-07, + 9.991350000000e-07, + 1.124700000000e-06,  \
+ 1.219100000000e-06, + 1.291100000000e-06, + 1.346900000000e-06, + 1.390900000000e-06, + 1.426100000000e-06,  \
+ 1.455100000000e-06, + 1.479400000000e-06, + 1.500500000000e-06, + 1.519200000000e-06, + 1.536100000000e-06,  \
+ 1.551700000000e-06, + 1.566200000000e-06, + 1.579900000000e-06, + 1.593000000000e-06, + 1.605500000000e-06,  \
+ 1.617700000000e-06, + 1.629400000000e-06, + 1.640900000000e-06, + 1.652100000000e-06, + 1.663200000000e-06,  \
+ 1.674000000000e-06, + 1.684700000000e-06, + 1.695200000000e-06, + 1.705700000000e-06, + 1.716000000000e-06,  \
+ 1.726300000000e-06, + 1.736400000000e-06, + 1.746500000000e-06, + 1.756500000000e-06, + 1.766500000000e-06,  \
+ 1.776400000000e-06, + 1.786300000000e-06, + 1.796200000000e-06, + 1.806000000000e-06, + 1.815800000000e-06,  \
+ 1.825500000000e-06, + 1.835200000000e-06, + 1.845000000000e-06, + 1.854600000000e-06, + 1.864300000000e-06,  \
+ 1.874000000000e-06, + 1.883600000000e-06, + 1.893300000000e-06, + 1.902900000000e-06, + 1.912500000000e-06,  \
+ 1.922200000000e-06, + 1.931800000000e-06, + 1.941400000000e-06, + 1.951000000000e-06, + 1.960600000000e-06,  \
+ 1.970300000000e-06, + 1.979900000000e-06, + 1.989500000000e-06, + 1.999200000000e-06, + 2.008800000000e-06,  \
+ 2.018400000000e-06, + 2.028100000000e-06, + 2.037700000000e-06, + 2.047400000000e-06, + 2.057100000000e-06,  \
+ 2.066800000000e-06, + 2.076500000000e-06, + 2.086200000000e-06, + 2.095900000000e-06, + 2.105600000000e-06,  \
+ 2.115300000000e-06, + 2.125100000000e-06, + 2.134900000000e-06, + 2.144600000000e-06, + 2.154400000000e-06,  \
+ 2.164200000000e-06, + 2.174000000000e-06, + 2.183900000000e-06, + 2.193700000000e-06, + 2.203600000000e-06 ]

.param id_pred_data_vg0.25=[ \
+ 3.354234286235e-07, + 6.017924533808e-07, + 8.126270950015e-07, + 9.789929754334e-07, + 1.109917866415e-06,  \
+ 1.212725073856e-06, + 1.293344266742e-06, + 1.356550783385e-06, + 1.406178034813e-06, + 1.445293219149e-06,  \
+ 1.476336756241e-06, + 1.501248407294e-06, + 1.521558533568e-06, + 1.538460728625e-06, + 1.552899539092e-06,  \
+ 1.565590500832e-06, + 1.577091024956e-06, + 1.587817969266e-06, + 1.598083727004e-06, + 1.608106504136e-06,  \
+ 1.618053802304e-06, + 1.628023101148e-06, + 1.638082421778e-06, + 1.648265133554e-06, + 1.658580572439e-06,  \
+ 1.669021075941e-06, + 1.679576357674e-06, + 1.690214030532e-06, + 1.700903885649e-06, + 1.711624599920e-06,  \
+ 1.722337697174e-06, + 1.733015960781e-06, + 1.743643033478e-06, + 1.754186014296e-06, + 1.764635339896e-06,  \
+ 1.774978827598e-06, + 1.785210256458e-06, + 1.795325661078e-06, + 1.805325314308e-06, + 1.815220639401e-06,  \
+ 1.825014128372e-06, + 1.834720515035e-06, + 1.844349048952e-06, + 1.853918092820e-06, + 1.863442980721e-06,  \
+ 1.872936609288e-06, + 1.882412593659e-06, + 1.891892025014e-06, + 1.901382443066e-06, + 1.910898845381e-06,  \
+ 1.920447425618e-06, + 1.930043299581e-06, + 1.939685489560e-06, + 1.949384418367e-06, + 1.959140058716e-06,  \
+ 1.968948854483e-06, + 1.978813390906e-06, + 1.988724061448e-06, + 1.998683012516e-06, + 2.008672072407e-06,  \
+ 2.018687241616e-06, + 2.028716098721e-06, + 2.038742525201e-06, + 2.048755559372e-06, + 2.058743120870e-06,  \
+ 2.068678340947e-06, + 2.078550949136e-06, + 2.088344035656e-06, + 2.098037498399e-06, + 2.107608634105e-06,  \
+ 2.117037788594e-06, + 2.126314157067e-06, + 2.135406680281e-06, + 2.144303321074e-06, + 2.152979448056e-06,  \
+ 2.161421634810e-06, + 2.169599997615e-06, + 2.177508363275e-06, + 2.185119585647e-06, + 2.192418833147e-06 ]

* Data table for Id-Vd at Vg = 0.26V
.param vd_data_vg0.26=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.26=[ \
+ 4.084390000000e-07, + 7.475790000000e-07, + 1.021900000000e-06, + 1.237500000000e-06, + 1.403200000000e-06,  \
+ 1.529600000000e-06, + 1.626600000000e-06, + 1.702100000000e-06, + 1.761600000000e-06, + 1.809200000000e-06,  \
+ 1.848100000000e-06, + 1.880600000000e-06, + 1.908400000000e-06, + 1.932900000000e-06, + 1.954800000000e-06,  \
+ 1.974800000000e-06, + 1.993300000000e-06, + 2.010600000000e-06, + 2.027100000000e-06, + 2.042800000000e-06,  \
+ 2.057800000000e-06, + 2.072400000000e-06, + 2.086600000000e-06, + 2.100500000000e-06, + 2.114000000000e-06,  \
+ 2.127300000000e-06, + 2.140300000000e-06, + 2.153200000000e-06, + 2.165900000000e-06, + 2.178400000000e-06,  \
+ 2.190800000000e-06, + 2.203100000000e-06, + 2.215300000000e-06, + 2.227400000000e-06, + 2.239400000000e-06,  \
+ 2.251400000000e-06, + 2.263300000000e-06, + 2.275100000000e-06, + 2.286800000000e-06, + 2.298600000000e-06,  \
+ 2.310200000000e-06, + 2.321900000000e-06, + 2.333500000000e-06, + 2.345000000000e-06, + 2.356600000000e-06,  \
+ 2.368100000000e-06, + 2.379600000000e-06, + 2.391000000000e-06, + 2.402500000000e-06, + 2.413900000000e-06,  \
+ 2.425300000000e-06, + 2.436800000000e-06, + 2.448200000000e-06, + 2.459600000000e-06, + 2.470900000000e-06,  \
+ 2.482300000000e-06, + 2.493700000000e-06, + 2.505100000000e-06, + 2.516500000000e-06, + 2.527800000000e-06,  \
+ 2.539200000000e-06, + 2.550600000000e-06, + 2.562000000000e-06, + 2.573400000000e-06, + 2.584700000000e-06,  \
+ 2.596100000000e-06, + 2.607500000000e-06, + 2.618900000000e-06, + 2.630400000000e-06, + 2.641800000000e-06,  \
+ 2.653200000000e-06, + 2.664600000000e-06, + 2.676100000000e-06, + 2.687500000000e-06, + 2.699000000000e-06,  \
+ 2.710500000000e-06, + 2.722000000000e-06, + 2.733500000000e-06, + 2.745000000000e-06, + 2.756500000000e-06 ]

.param id_pred_data_vg0.26=[ \
+ 4.076106051798e-07, + 7.359194569290e-07, + 9.995388973039e-07, + 1.210605914821e-06, + 1.379164314130e-06,  \
+ 1.513491224614e-06, + 1.620377115614e-06, + 1.705380127532e-06, + 1.773029871401e-06, + 1.826999141485e-06,  \
+ 1.870266150945e-06, + 1.905216195155e-06, + 1.933775956786e-06, + 1.957473814400e-06, + 1.977528609132e-06,  \
+ 1.994895574171e-06, + 2.010320349655e-06, + 2.024387595156e-06, + 2.037540180027e-06, + 2.050108014373e-06,  \
+ 2.062333087451e-06, + 2.074400581478e-06, + 2.086425811285e-06, + 2.098482800648e-06, + 2.110621380780e-06,  \
+ 2.122862297256e-06, + 2.135198319593e-06, + 2.147627710656e-06, + 2.160124513466e-06, + 2.172666108891e-06,  \
+ 2.185224689129e-06, + 2.197772701038e-06, + 2.210284210378e-06, + 2.222743423772e-06, + 2.235124588879e-06,  \
+ 2.247411212011e-06, + 2.259598577439e-06, + 2.271680432386e-06, + 2.283658182023e-06, + 2.295529338880e-06,  \
+ 2.307302338522e-06, + 2.318989909327e-06, + 2.330601946596e-06, + 2.342153256905e-06, + 2.353650074838e-06,  \
+ 2.365122199990e-06, + 2.376574002483e-06, + 2.388022548985e-06, + 2.399484346824e-06, + 2.410967454125e-06,  \
+ 2.422485513307e-06, + 2.434039633954e-06, + 2.445644554427e-06, + 2.457296932334e-06, + 2.469008177286e-06,  \
+ 2.480763832864e-06, + 2.492567568879e-06, + 2.504413514544e-06, + 2.516292265682e-06, + 2.528188269935e-06,  \
+ 2.540088867136e-06, + 2.551987463448e-06, + 2.563861453382e-06, + 2.575691905804e-06, + 2.587468338788e-06,  \
+ 2.599156960059e-06, + 2.610741798890e-06, + 2.622201936902e-06, + 2.633514509398e-06, + 2.644653204698e-06,  \
+ 2.655590662926e-06, + 2.666314012458e-06, + 2.676786250504e-06, + 2.686984944376e-06, + 2.696897297483e-06,  \
+ 2.706483619477e-06, + 2.715732041452e-06, + 2.724609794313e-06, + 2.733109020028e-06, + 2.741195385170e-06 ]

* Data table for Id-Vd at Vg = 0.27V
.param vd_data_vg0.27=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.27=[ \
+ 4.811210000000e-07, + 8.890820000000e-07, + 1.226700000000e-06, + 1.498600000000e-06, + 1.712200000000e-06,  \
+ 1.877800000000e-06, + 2.006400000000e-06, + 2.106900000000e-06, + 2.186400000000e-06, + 2.249900000000e-06,  \
+ 2.301600000000e-06, + 2.344500000000e-06, + 2.381000000000e-06, + 2.412700000000e-06, + 2.440800000000e-06,  \
+ 2.466200000000e-06, + 2.489600000000e-06, + 2.511300000000e-06, + 2.531700000000e-06, + 2.551100000000e-06,  \
+ 2.569700000000e-06, + 2.587500000000e-06, + 2.604800000000e-06, + 2.621600000000e-06, + 2.638000000000e-06,  \
+ 2.654000000000e-06, + 2.669700000000e-06, + 2.685100000000e-06, + 2.700300000000e-06, + 2.715300000000e-06,  \
+ 2.730100000000e-06, + 2.744800000000e-06, + 2.759200000000e-06, + 2.773600000000e-06, + 2.787800000000e-06,  \
+ 2.802000000000e-06, + 2.816000000000e-06, + 2.830000000000e-06, + 2.843800000000e-06, + 2.857600000000e-06,  \
+ 2.871300000000e-06, + 2.885000000000e-06, + 2.898600000000e-06, + 2.912200000000e-06, + 2.925700000000e-06,  \
+ 2.939200000000e-06, + 2.952700000000e-06, + 2.966100000000e-06, + 2.979500000000e-06, + 2.992800000000e-06,  \
+ 3.006100000000e-06, + 3.019400000000e-06, + 3.032700000000e-06, + 3.046000000000e-06, + 3.059200000000e-06,  \
+ 3.072500000000e-06, + 3.085700000000e-06, + 3.098900000000e-06, + 3.112100000000e-06, + 3.125300000000e-06,  \
+ 3.138500000000e-06, + 3.151700000000e-06, + 3.164900000000e-06, + 3.178100000000e-06, + 3.191200000000e-06,  \
+ 3.204400000000e-06, + 3.217600000000e-06, + 3.230800000000e-06, + 3.243900000000e-06, + 3.257100000000e-06,  \
+ 3.270300000000e-06, + 3.283500000000e-06, + 3.296700000000e-06, + 3.309900000000e-06, + 3.323100000000e-06,  \
+ 3.336300000000e-06, + 3.349500000000e-06, + 3.362700000000e-06, + 3.375900000000e-06, + 3.389200000000e-06 ]

.param id_pred_data_vg0.27=[ \
+ 4.852415804635e-07, + 8.815071487334e-07, + 1.204168656841e-06, + 1.466180547141e-06, + 1.678416447248e-06,  \
+ 1.849984037108e-06, + 1.988452131627e-06, + 2.100105484715e-06, + 2.190153481934e-06, + 2.262871385028e-06,  \
+ 2.321784213564e-06, + 2.369764188188e-06, + 2.409151311440e-06, + 2.441851247568e-06, + 2.469389710313e-06,  \
+ 2.493001229595e-06, + 2.513655417715e-06, + 2.532133494242e-06, + 2.549044147599e-06, + 2.564862552390e-06,  \
+ 2.579935498943e-06, + 2.594536908873e-06, + 2.608868371681e-06, + 2.623063555802e-06, + 2.637225179569e-06,  \
+ 2.651405138749e-06, + 2.665640186024e-06, + 2.679942954273e-06, + 2.694306513149e-06, + 2.708727151912e-06,  \
+ 2.723176421568e-06, + 2.737641043495e-06, + 2.752097061602e-06, + 2.766517809505e-06, + 2.780893601084e-06,  \
+ 2.795201980916e-06, + 2.809432617141e-06, + 2.823579061442e-06, + 2.837641382030e-06, + 2.851611498045e-06,  \
+ 2.865495866899e-06, + 2.879305238821e-06, + 2.893046948884e-06, + 2.906731515395e-06, + 2.920372935478e-06,  \
+ 2.933986197604e-06, + 2.947588041025e-06, + 2.961185600725e-06, + 2.974794192596e-06, + 2.988426103911e-06,  \
+ 3.002090325026e-06, + 3.015793354280e-06, + 3.029533522749e-06, + 3.043329234060e-06, + 3.057165554310e-06,  \
+ 3.071050814469e-06, + 3.084962900175e-06, + 3.098905908701e-06, + 3.112871204394e-06, + 3.126826959488e-06,  \
+ 3.140778558191e-06, + 3.154693549732e-06, + 3.168553066644e-06, + 3.182339132763e-06, + 3.196023294549e-06,  \
+ 3.209585374861e-06, + 3.222996801924e-06, + 3.236224620196e-06, + 3.249246865380e-06, + 3.262031395934e-06,  \
+ 3.274548007539e-06, + 3.286773753644e-06, + 3.298672781966e-06, + 3.310214833618e-06, + 3.321368012621e-06,  \
+ 3.332112701173e-06, + 3.342421550769e-06, + 3.352254152560e-06, + 3.361595513525e-06, + 3.370409831405e-06 ]

* Data table for Id-Vd at Vg = 0.28V
.param vd_data_vg0.28=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.28=[ \
+ 5.560310000000e-07, + 1.036400000000e-06, + 1.442300000000e-06, + 1.776700000000e-06, + 2.045400000000e-06,  \
+ 2.257800000000e-06, + 2.424700000000e-06, + 2.556400000000e-06, + 2.661000000000e-06, + 2.744700000000e-06,  \
+ 2.812600000000e-06, + 2.868800000000e-06, + 2.916100000000e-06, + 2.956900000000e-06, + 2.992700000000e-06,  \
+ 3.024800000000e-06, + 3.054000000000e-06, + 3.080900000000e-06, + 3.106100000000e-06, + 3.129800000000e-06,  \
+ 3.152400000000e-06, + 3.174000000000e-06, + 3.194800000000e-06, + 3.214900000000e-06, + 3.234500000000e-06,  \
+ 3.253600000000e-06, + 3.272200000000e-06, + 3.290500000000e-06, + 3.308400000000e-06, + 3.326100000000e-06,  \
+ 3.343500000000e-06, + 3.360600000000e-06, + 3.377600000000e-06, + 3.394400000000e-06, + 3.411000000000e-06,  \
+ 3.427500000000e-06, + 3.443800000000e-06, + 3.460100000000e-06, + 3.476200000000e-06, + 3.492200000000e-06,  \
+ 3.508100000000e-06, + 3.523900000000e-06, + 3.539700000000e-06, + 3.555300000000e-06, + 3.571000000000e-06,  \
+ 3.586500000000e-06, + 3.602000000000e-06, + 3.617400000000e-06, + 3.632800000000e-06, + 3.648200000000e-06,  \
+ 3.663500000000e-06, + 3.678800000000e-06, + 3.694000000000e-06, + 3.709200000000e-06, + 3.724400000000e-06,  \
+ 3.739600000000e-06, + 3.754700000000e-06, + 3.769800000000e-06, + 3.784900000000e-06, + 3.800000000000e-06,  \
+ 3.815100000000e-06, + 3.830100000000e-06, + 3.845100000000e-06, + 3.860200000000e-06, + 3.875200000000e-06,  \
+ 3.890200000000e-06, + 3.905200000000e-06, + 3.920200000000e-06, + 3.935100000000e-06, + 3.950100000000e-06,  \
+ 3.965100000000e-06, + 3.980100000000e-06, + 3.995000000000e-06, + 4.010000000000e-06, + 4.025000000000e-06,  \
+ 4.040000000000e-06, + 4.054900000000e-06, + 4.069900000000e-06, + 4.084900000000e-06, + 4.099900000000e-06 ]

.param id_pred_data_vg0.28=[ \
+ 5.667030200129e-07, + 1.035695968312e-06, + 1.422750356141e-06, + 1.741349988151e-06, + 2.002974542847e-06,  \
+ 2.217367655248e-06, + 2.392755377514e-06, + 2.536080137361e-06, + 2.653153278516e-06, + 2.748838232947e-06,  \
+ 2.827183998306e-06, + 2.891561016440e-06, + 2.944735952042e-06, + 2.989009772136e-06, + 3.026255035365e-06,  \
+ 3.058001166210e-06, + 3.085495354753e-06, + 3.109730605502e-06, + 3.131511111860e-06, + 3.151478813379e-06,  \
+ 3.170138315909e-06, + 3.187864131178e-06, + 3.204965378245e-06, + 3.221657389076e-06, + 3.238109002268e-06,  \
+ 3.254436305724e-06, + 3.270717170381e-06, + 3.286999963166e-06, + 3.303302974018e-06, + 3.319650295452e-06,  \
+ 3.336031622894e-06, + 3.352437051944e-06, + 3.368863990545e-06, + 3.385282816453e-06, + 3.401683261472e-06,  \
+ 3.418057603994e-06, + 3.434388145251e-06, + 3.450661079114e-06, + 3.466871085038e-06, + 3.483028558549e-06,  \
+ 3.499116292005e-06, + 3.515150820022e-06, + 3.531142601787e-06, + 3.547084415914e-06, + 3.563003792806e-06,  \
+ 3.578902724257e-06, + 3.594791287469e-06, + 3.610692729126e-06, + 3.626601387623e-06, + 3.642535830295e-06,  \
+ 3.658503478619e-06, + 3.674508625409e-06, + 3.690556559377e-06, + 3.706644565682e-06, + 3.722772316905e-06,  \
+ 3.738928426174e-06, + 3.755106549761e-06, + 3.771301580855e-06, + 3.787491373259e-06, + 3.803659092227e-06,  \
+ 3.819785429187e-06, + 3.835848965537e-06, + 3.851822812067e-06, + 3.867681662086e-06, + 3.883390877490e-06,  \
+ 3.898932327502e-06, + 3.914257345059e-06, + 3.929351278202e-06, + 3.944162081098e-06, + 3.958669185522e-06,  \
+ 3.972827721554e-06, + 3.986607334809e-06, + 3.999968298558e-06, + 4.012888721263e-06, + 4.025315206491e-06,  \
+ 4.037220041937e-06, + 4.048575165143e-06, + 4.059347002112e-06, + 4.069505625921e-06, + 4.079005157109e-06 ]

* Data table for Id-Vd at Vg = 0.29V
.param vd_data_vg0.29=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.29=[ \
+ 6.319470000000e-07, + 1.186900000000e-06, + 1.664600000000e-06, + 2.066400000000e-06, + 2.396300000000e-06,  \
+ 2.662200000000e-06, + 2.874400000000e-06, + 3.043600000000e-06, + 3.179000000000e-06, + 3.287800000000e-06,  \
+ 3.376100000000e-06, + 3.448800000000e-06, + 3.509700000000e-06, + 3.561700000000e-06, + 3.607000000000e-06,  \
+ 3.647200000000e-06, + 3.683500000000e-06, + 3.716700000000e-06, + 3.747400000000e-06, + 3.776200000000e-06,  \
+ 3.803400000000e-06, + 3.829300000000e-06, + 3.854100000000e-06, + 3.878000000000e-06, + 3.901100000000e-06,  \
+ 3.923600000000e-06, + 3.945500000000e-06, + 3.966800000000e-06, + 3.987800000000e-06, + 4.008300000000e-06,  \
+ 4.028500000000e-06, + 4.048500000000e-06, + 4.068100000000e-06, + 4.087500000000e-06, + 4.106600000000e-06,  \
+ 4.125600000000e-06, + 4.144400000000e-06, + 4.163000000000e-06, + 4.181500000000e-06, + 4.199800000000e-06,  \
+ 4.218000000000e-06, + 4.236100000000e-06, + 4.254100000000e-06, + 4.271900000000e-06, + 4.289700000000e-06,  \
+ 4.307400000000e-06, + 4.325000000000e-06, + 4.342600000000e-06, + 4.360100000000e-06, + 4.377500000000e-06,  \
+ 4.394900000000e-06, + 4.412200000000e-06, + 4.429400000000e-06, + 4.446600000000e-06, + 4.463800000000e-06,  \
+ 4.480900000000e-06, + 4.498000000000e-06, + 4.515100000000e-06, + 4.532100000000e-06, + 4.549100000000e-06,  \
+ 4.566000000000e-06, + 4.583000000000e-06, + 4.599900000000e-06, + 4.616800000000e-06, + 4.633700000000e-06,  \
+ 4.650500000000e-06, + 4.667400000000e-06, + 4.684200000000e-06, + 4.701000000000e-06, + 4.717800000000e-06,  \
+ 4.734600000000e-06, + 4.751400000000e-06, + 4.768100000000e-06, + 4.784900000000e-06, + 4.801700000000e-06,  \
+ 4.818400000000e-06, + 4.835200000000e-06, + 4.851900000000e-06, + 4.868600000000e-06, + 4.885400000000e-06 ]

.param id_pred_data_vg0.29=[ \
+ 6.503488111775e-07, + 1.195480508613e-06, + 1.651201637287e-06, + 2.031215262832e-06, + 2.347348890908e-06,  \
+ 2.609791554278e-06, + 2.827268253895e-06, + 3.007243794855e-06, + 3.156062557537e-06, + 3.279096927145e-06,  \
+ 3.380906236998e-06, + 3.465326080914e-06, + 3.535564155754e-06, + 3.594307345338e-06, + 3.643800482678e-06,  \
+ 3.685896517709e-06, + 3.722119527083e-06, + 3.753720739041e-06, + 3.781742470892e-06, + 3.807003304246e-06,  \
+ 3.830179957731e-06, + 3.851798101095e-06, + 3.872272936860e-06, + 3.891950327670e-06, + 3.911078692909e-06,  \
+ 3.929843423975e-06, + 3.948381026930e-06, + 3.966792537540e-06, + 3.985155790360e-06, + 4.003502817795e-06,  \
+ 4.021869835924e-06, + 4.040256899316e-06, + 4.058671947860e-06, + 4.077103603777e-06, + 4.095558324479e-06,  \
+ 4.114017174288e-06, + 4.132466610827e-06, + 4.150895347266e-06, + 4.169316971456e-06, + 4.187705781078e-06,  \
+ 4.206065532344e-06, + 4.224405092828e-06, + 4.242716831868e-06, + 4.261017384124e-06, + 4.279308632249e-06,  \
+ 4.297596278775e-06, + 4.315897458582e-06, + 4.334207478678e-06, + 4.352544419817e-06, + 4.370917849883e-06,  \
+ 4.389316472952e-06, + 4.407762353367e-06, + 4.426235536812e-06, + 4.444746773515e-06, + 4.463298091650e-06,  \
+ 4.481860014494e-06, + 4.500437562456e-06, + 4.519002031884e-06, + 4.537545155472e-06, + 4.556041039905e-06,  \
+ 4.574458407660e-06, + 4.592784553097e-06, + 4.610977962329e-06, + 4.629017785192e-06, + 4.646852880796e-06,  \
+ 4.664457901526e-06, + 4.681795621764e-06, + 4.698823286162e-06, + 4.715500185739e-06, + 4.731788249046e-06,  \
+ 4.747647790282e-06, + 4.763038086821e-06, + 4.777902713613e-06, + 4.792225327037e-06, + 4.805951220987e-06,  \
+ 4.819043715543e-06, + 4.831445389755e-06, + 4.843145425184e-06, + 4.854108155996e-06, + 4.864265429205e-06 ]

* Data table for Id-Vd at Vg = 0.30V
.param vd_data_vg0.30=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.30=[ \
+ 7.078840000000e-07, + 1.338300000000e-06, + 1.890000000000e-06, + 2.362500000000e-06, + 2.758300000000e-06,  \
+ 3.083600000000e-06, + 3.347500000000e-06, + 3.560600000000e-06, + 3.732700000000e-06, + 3.871800000000e-06,  \
+ 3.985000000000e-06, + 4.078200000000e-06, + 4.155800000000e-06, + 4.221800000000e-06, + 4.278700000000e-06,  \
+ 4.328800000000e-06, + 4.373600000000e-06, + 4.414200000000e-06, + 4.451500000000e-06, + 4.486200000000e-06,  \
+ 4.518800000000e-06, + 4.549600000000e-06, + 4.578900000000e-06, + 4.607100000000e-06, + 4.634200000000e-06,  \
+ 4.660400000000e-06, + 4.685800000000e-06, + 4.710600000000e-06, + 4.734800000000e-06, + 4.758500000000e-06,  \
+ 4.781700000000e-06, + 4.804500000000e-06, + 4.827000000000e-06, + 4.849200000000e-06, + 4.871000000000e-06,  \
+ 4.892600000000e-06, + 4.914000000000e-06, + 4.935100000000e-06, + 4.956100000000e-06, + 4.976800000000e-06,  \
+ 4.997400000000e-06, + 5.017800000000e-06, + 5.038100000000e-06, + 5.058300000000e-06, + 5.078300000000e-06,  \
+ 5.098200000000e-06, + 5.118000000000e-06, + 5.137800000000e-06, + 5.157400000000e-06, + 5.176900000000e-06,  \
+ 5.196400000000e-06, + 5.215700000000e-06, + 5.235000000000e-06, + 5.254300000000e-06, + 5.273500000000e-06,  \
+ 5.292600000000e-06, + 5.311700000000e-06, + 5.330700000000e-06, + 5.349700000000e-06, + 5.368600000000e-06,  \
+ 5.387500000000e-06, + 5.406400000000e-06, + 5.425200000000e-06, + 5.444000000000e-06, + 5.462700000000e-06,  \
+ 5.481400000000e-06, + 5.500100000000e-06, + 5.518800000000e-06, + 5.537500000000e-06, + 5.556100000000e-06,  \
+ 5.574700000000e-06, + 5.593300000000e-06, + 5.611800000000e-06, + 5.630400000000e-06, + 5.648900000000e-06,  \
+ 5.667400000000e-06, + 5.686000000000e-06, + 5.704500000000e-06, + 5.722900000000e-06, + 5.741400000000e-06 ]

.param id_pred_data_vg0.30=[ \
+ 7.346443453571e-07, + 1.357968139928e-06, + 1.885468955152e-06, + 2.330768329557e-06, + 2.705799488467e-06,  \
+ 3.020970834768e-06, + 3.285329657956e-06, + 3.506719367579e-06, + 3.691908787005e-06, + 3.846712206723e-06,  \
+ 3.976120096922e-06, + 4.084414104000e-06, + 4.175199719612e-06, + 4.251566970197e-06, + 4.316111790104e-06,  \
+ 4.371028626338e-06, + 4.418149837875e-06, + 4.459014344320e-06, + 4.494872064242e-06, + 4.526795964921e-06,  \
+ 4.555631276162e-06, + 4.582100336847e-06, + 4.606746897480e-06, + 4.630041948985e-06, + 4.652349616663e-06,  \
+ 4.673944204114e-06, + 4.695056104538e-06, + 4.715838222182e-06, + 4.736422451970e-06, + 4.756912312587e-06,  \
+ 4.777345802722e-06, + 4.797777510248e-06, + 4.818220368179e-06, + 4.838707609451e-06, + 4.859228602072e-06,  \
+ 4.879779335170e-06, + 4.900373214696e-06, + 4.920991505060e-06, + 4.941638626406e-06, + 4.962293314748e-06,  \
+ 4.982969840057e-06, + 5.003656715417e-06, + 5.024359006711e-06, + 5.045078687544e-06, + 5.065807408755e-06,  \
+ 5.086573492008e-06, + 5.107362676426e-06, + 5.128184129717e-06, + 5.149050048203e-06, + 5.169938049221e-06,  \
+ 5.190883275645e-06, + 5.211862553551e-06, + 5.232877365415e-06, + 5.253919989627e-06, + 5.274988461679e-06,  \
+ 5.296062372508e-06, + 5.317127206581e-06, + 5.338169648894e-06, + 5.359169017538e-06, + 5.380085531215e-06,  \
+ 5.400891204772e-06, + 5.421566638688e-06, + 5.442072679216e-06, + 5.462353001349e-06, + 5.482394954015e-06,  \
+ 5.502142412297e-06, + 5.521566690732e-06, + 5.540602433030e-06, + 5.559211904256e-06, + 5.577334104601e-06,  \
+ 5.594944886980e-06, + 5.611984088318e-06, + 5.628408453049e-06, + 5.644160919474e-06, + 5.659220505549e-06,  \
+ 5.673495525116e-06, + 5.686984427484e-06, + 5.699619996449e-06, + 5.711372314181e-06, + 5.722182322643e-06 ]

* Data table for Id-Vd at Vg = 0.31V
.param vd_data_vg0.31=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.31=[ \
+ 7.830880000000e-07, + 1.489100000000e-06, + 2.115400000000e-06, + 2.660700000000e-06, + 3.125800000000e-06,  \
+ 3.514900000000e-06, + 3.836000000000e-06, + 4.099000000000e-06, + 4.313500000000e-06, + 4.488500000000e-06,  \
+ 4.631600000000e-06, + 4.749500000000e-06, + 4.847600000000e-06, + 4.930400000000e-06, + 5.001500000000e-06,  \
+ 5.063600000000e-06, + 5.118600000000e-06, + 5.168100000000e-06, + 5.213200000000e-06, + 5.254800000000e-06,  \
+ 5.293500000000e-06, + 5.329900000000e-06, + 5.364500000000e-06, + 5.397400000000e-06, + 5.428900000000e-06,  \
+ 5.459300000000e-06, + 5.488600000000e-06, + 5.517100000000e-06, + 5.544900000000e-06, + 5.572000000000e-06,  \
+ 5.598500000000e-06, + 5.624400000000e-06, + 5.650000000000e-06, + 5.675000000000e-06, + 5.699800000000e-06,  \
+ 5.724100000000e-06, + 5.748200000000e-06, + 5.772000000000e-06, + 5.795500000000e-06, + 5.818800000000e-06,  \
+ 5.841800000000e-06, + 5.864700000000e-06, + 5.887400000000e-06, + 5.909900000000e-06, + 5.932200000000e-06,  \
+ 5.954400000000e-06, + 5.976500000000e-06, + 5.998400000000e-06, + 6.020200000000e-06, + 6.041900000000e-06,  \
+ 6.063500000000e-06, + 6.085000000000e-06, + 6.106400000000e-06, + 6.127700000000e-06, + 6.148900000000e-06,  \
+ 6.170000000000e-06, + 6.191100000000e-06, + 6.212100000000e-06, + 6.233100000000e-06, + 6.254000000000e-06,  \
+ 6.274800000000e-06, + 6.295600000000e-06, + 6.316300000000e-06, + 6.337000000000e-06, + 6.357600000000e-06,  \
+ 6.378200000000e-06, + 6.398800000000e-06, + 6.419300000000e-06, + 6.439800000000e-06, + 6.460200000000e-06,  \
+ 6.480600000000e-06, + 6.501000000000e-06, + 6.521400000000e-06, + 6.541700000000e-06, + 6.562000000000e-06,  \
+ 6.582300000000e-06, + 6.602500000000e-06, + 6.622800000000e-06, + 6.643000000000e-06, + 6.663200000000e-06 ]

.param id_pred_data_vg0.31=[ \
+ 8.182539022528e-07, + 1.520556397736e-06, + 2.121807192452e-06, + 2.635279379319e-06, + 3.072764229728e-06,  \
+ 3.444665344432e-06, + 3.760185027204e-06, + 4.027392715216e-06, + 4.253350271028e-06, + 4.444202204468e-06,  \
+ 4.605325448210e-06, + 4.741357115563e-06, + 4.856294617639e-06, + 4.953591997037e-06, + 5.036199945607e-06,  \
+ 5.106644821353e-06, + 5.167064664420e-06, + 5.219289305387e-06, + 5.264839655865e-06, + 5.305013837642e-06,  \
+ 5.340884308680e-06, + 5.373334824981e-06, + 5.403123777796e-06, + 5.430844612420e-06, + 5.456989583763e-06,  \
+ 5.481953230628e-06, + 5.506058278115e-06, + 5.529550107894e-06, + 5.552626535064e-06, + 5.575444993156e-06,  \
+ 5.598086863756e-06, + 5.620672018267e-06, + 5.643238055200e-06, + 5.665817589033e-06, + 5.688446708518e-06,  \
+ 5.711142657674e-06, + 5.733894140576e-06, + 5.756712744187e-06, + 5.779609055026e-06, + 5.802559826407e-06,  \
+ 5.825570779052e-06, + 5.848651107954e-06, + 5.871774646948e-06, + 5.894954410905e-06, + 5.918198667132e-06,  \
+ 5.941483759671e-06, + 5.964828533251e-06, + 5.988220655126e-06, + 6.011662862875e-06, + 6.035169008101e-06,  \
+ 6.058712733648e-06, + 6.082311592763e-06, + 6.105933589424e-06, + 6.129586909083e-06, + 6.153245385576e-06,  \
+ 6.176908864290e-06, + 6.200542693477e-06, + 6.224125972949e-06, + 6.247644887480e-06, + 6.271054007811e-06,  \
+ 6.294315107880e-06, + 6.317398238025e-06, + 6.340270711007e-06, + 6.362878484651e-06, + 6.385189590219e-06,  \
+ 6.407131204469e-06, + 6.428665801650e-06, + 6.449764259742e-06, + 6.470341149907e-06, + 6.490362557088e-06,  \
+ 6.509769727927e-06, + 6.528505909955e-06, + 6.546513668582e-06, + 6.563752122020e-06, + 6.580154831681e-06,  \
+ 6.595664381166e-06, + 6.610242480747e-06, + 6.623836798099e-06, + 6.636399721174e-06, + 6.647882401012e-06 ]

* Data table for Id-Vd at Vg = 0.32V
.param vd_data_vg0.32=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.32=[ \
+ 8.570000000000e-07, + 1.637700000000e-06, + 2.338800000000e-06, + 2.957700000000e-06, + 3.494000000000e-06,  \
+ 3.950300000000e-06, + 4.332900000000e-06, + 4.650600000000e-06, + 4.913100000000e-06, + 5.129300000000e-06,  \
+ 5.307400000000e-06, + 5.454600000000e-06, + 5.577100000000e-06, + 5.680400000000e-06, + 5.768500000000e-06,  \
+ 5.844900000000e-06, + 5.912100000000e-06, + 5.972100000000e-06, + 6.026400000000e-06, + 6.076100000000e-06,  \
+ 6.122000000000e-06, + 6.164900000000e-06, + 6.205300000000e-06, + 6.243600000000e-06, + 6.280100000000e-06,  \
+ 6.315100000000e-06, + 6.348800000000e-06, + 6.381400000000e-06, + 6.413000000000e-06, + 6.443800000000e-06,  \
+ 6.473800000000e-06, + 6.503200000000e-06, + 6.531900000000e-06, + 6.560100000000e-06, + 6.587900000000e-06,  \
+ 6.615200000000e-06, + 6.642100000000e-06, + 6.668600000000e-06, + 6.694800000000e-06, + 6.720700000000e-06,  \
+ 6.746400000000e-06, + 6.771700000000e-06, + 6.796900000000e-06, + 6.821800000000e-06, + 6.846500000000e-06,  \
+ 6.871000000000e-06, + 6.895400000000e-06, + 6.919600000000e-06, + 6.943600000000e-06, + 6.967500000000e-06,  \
+ 6.991300000000e-06, + 7.014900000000e-06, + 7.038400000000e-06, + 7.061800000000e-06, + 7.085100000000e-06,  \
+ 7.108300000000e-06, + 7.131400000000e-06, + 7.154400000000e-06, + 7.177300000000e-06, + 7.200200000000e-06,  \
+ 7.222900000000e-06, + 7.245700000000e-06, + 7.268300000000e-06, + 7.290900000000e-06, + 7.313400000000e-06,  \
+ 7.335800000000e-06, + 7.358200000000e-06, + 7.380600000000e-06, + 7.402900000000e-06, + 7.425100000000e-06,  \
+ 7.447400000000e-06, + 7.469500000000e-06, + 7.491700000000e-06, + 7.513800000000e-06, + 7.535800000000e-06,  \
+ 7.557800000000e-06, + 7.579800000000e-06, + 7.601800000000e-06, + 7.623700000000e-06, + 7.645600000000e-06 ]

.param id_pred_data_vg0.32=[ \
+ 9.000972931972e-07, + 1.681071589701e-06, + 2.356989207328e-06, + 2.940545382444e-06, + 3.443157766014e-06,  \
+ 3.875065594912e-06, + 4.245406271366e-06, + 4.562345857266e-06, + 4.833094753849e-06, + 5.064051947556e-06,  \
+ 5.260851685307e-06, + 5.428439180832e-06, + 5.571147303272e-06, + 5.692753111362e-06, + 5.796542245662e-06,  \
+ 5.885363207199e-06, + 5.961656206637e-06, + 6.027547715348e-06, + 6.084828128223e-06, + 6.135043076938e-06,  \
+ 6.179495685501e-06, + 6.219300812518e-06, + 6.255366115511e-06, + 6.288478762144e-06, + 6.319277417788e-06,  \
+ 6.348288661684e-06, + 6.375947086781e-06, + 6.402600993169e-06, + 6.428529632103e-06, + 6.453957394115e-06,  \
+ 6.479054409283e-06, + 6.503959302790e-06, + 6.528770409204e-06, + 6.553554849233e-06, + 6.578374450328e-06,  \
+ 6.603247602470e-06, + 6.628219271079e-06, + 6.653283453488e-06, + 6.678459631075e-06, + 6.703732651658e-06,  \
+ 6.729110609740e-06, + 6.754605019523e-06, + 6.780190979043e-06, + 6.805872835685e-06, + 6.831634163973e-06,  \
+ 6.857493262942e-06, + 6.883425803608e-06, + 6.909438525327e-06, + 6.935527926544e-06, + 6.961670806049e-06,  \
+ 6.987875131017e-06, + 7.014123293629e-06, + 7.040404088912e-06, + 7.066713478707e-06, + 7.093028625604e-06,  \
+ 7.119314977899e-06, + 7.145559520723e-06, + 7.171738361649e-06, + 7.197815484687e-06, + 7.223744069051e-06,  \
+ 7.249508971654e-06, + 7.275040279637e-06, + 7.300307788682e-06, + 7.325269980356e-06, + 7.349868656092e-06,  \
+ 7.374056694971e-06, + 7.397761346510e-06, + 7.420929432556e-06, + 7.443510748999e-06, + 7.465454473277e-06,  \
+ 7.486684526157e-06, + 7.507144182455e-06, + 7.526774788857e-06, + 7.545515454694e-06, + 7.563289045720e-06,  \
+ 7.580060300825e-06, + 7.595757124363e-06, + 7.610347238369e-06, + 7.623741266798e-06, + 7.635905785719e-06 ]

* Data table for Id-Vd at Vg = 0.33V
.param vd_data_vg0.33=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.33=[ \
+ 9.292130000000e-07, + 1.783400000000e-06, + 2.558400000000e-06, + 3.250900000000e-06, + 3.859200000000e-06,  \
+ 4.384600000000e-06, + 4.831800000000e-06, + 5.208500000000e-06, + 5.523500000000e-06, + 5.785900000000e-06,  \
+ 6.003900000000e-06, + 6.185100000000e-06, + 6.336400000000e-06, + 6.463700000000e-06, + 6.572200000000e-06,  \
+ 6.665700000000e-06, + 6.747400000000e-06, + 6.819900000000e-06, + 6.884900000000e-06, + 6.944000000000e-06,  \
+ 6.998300000000e-06, + 7.048700000000e-06, + 7.095800000000e-06, + 7.140200000000e-06, + 7.182300000000e-06,  \
+ 7.222500000000e-06, + 7.261000000000e-06, + 7.298100000000e-06, + 7.333900000000e-06, + 7.368700000000e-06,  \
+ 7.402500000000e-06, + 7.435500000000e-06, + 7.467700000000e-06, + 7.499300000000e-06, + 7.530200000000e-06,  \
+ 7.560600000000e-06, + 7.590500000000e-06, + 7.619900000000e-06, + 7.648900000000e-06, + 7.677600000000e-06,  \
+ 7.705900000000e-06, + 7.733900000000e-06, + 7.761600000000e-06, + 7.789000000000e-06, + 7.816200000000e-06,  \
+ 7.843100000000e-06, + 7.869800000000e-06, + 7.896300000000e-06, + 7.922600000000e-06, + 7.948700000000e-06,  \
+ 7.974700000000e-06, + 8.000500000000e-06, + 8.026100000000e-06, + 8.051600000000e-06, + 8.077000000000e-06,  \
+ 8.102300000000e-06, + 8.127400000000e-06, + 8.152400000000e-06, + 8.177300000000e-06, + 8.202200000000e-06,  \
+ 8.226900000000e-06, + 8.251500000000e-06, + 8.276100000000e-06, + 8.300500000000e-06, + 8.324900000000e-06,  \
+ 8.349200000000e-06, + 8.373500000000e-06, + 8.397600000000e-06, + 8.421800000000e-06, + 8.445800000000e-06,  \
+ 8.469800000000e-06, + 8.493800000000e-06, + 8.517600000000e-06, + 8.541500000000e-06, + 8.565300000000e-06,  \
+ 8.589000000000e-06, + 8.612700000000e-06, + 8.636400000000e-06, + 8.660000000000e-06, + 8.683600000000e-06 ]

.param id_pred_data_vg0.33=[ \
+ 9.793627395993e-07, + 1.837807503762e-06, + 2.588389324956e-06, + 3.243032260798e-06, + 3.812617069343e-06,  \
+ 4.307022609282e-06, + 4.735198890558e-06, + 5.105215823278e-06, + 5.424353548733e-06, + 5.699104804080e-06,  \
+ 5.935293520452e-06, + 6.138083408587e-06, + 6.312094301393e-06, + 6.461373632192e-06, + 6.589511758648e-06,  \
+ 6.699620280415e-06, + 6.794479486416e-06, + 6.876484549139e-06, + 6.947693764232e-06, + 7.009915134404e-06,  \
+ 7.064686651574e-06, + 7.113347746781e-06, + 7.157013060350e-06, + 7.196648803074e-06, + 7.233074484247e-06,  \
+ 7.266953180078e-06, + 7.298851105588e-06, + 7.329243744607e-06, + 7.358504299191e-06, + 7.386927063635e-06,  \
+ 7.414796218654e-06, + 7.442276109941e-06, + 7.469533884432e-06, + 7.496681682824e-06, + 7.523817112087e-06,  \
+ 7.550990703749e-06, + 7.578230579384e-06, + 7.605618011439e-06, + 7.633116329089e-06, + 7.660759729333e-06,  \
+ 7.688558634982e-06, + 7.716495310888e-06, + 7.744580634608e-06, + 7.772780518280e-06, + 7.801115862094e-06,  \
+ 7.829569040041e-06, + 7.858128810767e-06, + 7.886785897426e-06, + 7.915539845271e-06, + 7.944368917379e-06,  \
+ 7.973245938047e-06, + 8.002188042155e-06, + 8.031151846808e-06, + 8.060148757068e-06, + 8.089121865851e-06,  \
+ 8.118061741698e-06, + 8.146931359079e-06, + 8.175710645446e-06, + 8.204358255171e-06, + 8.232837899413e-06,  \
+ 8.261082439276e-06, + 8.289092984342e-06, + 8.316772100443e-06, + 8.344087982550e-06, + 8.370982732231e-06,  \
+ 8.397409637837e-06, + 8.423287417827e-06, + 8.448554726783e-06, + 8.473148673147e-06, + 8.497000999341e-06,  \
+ 8.520075853085e-06, + 8.542267969460e-06, + 8.563535120629e-06, + 8.583784710936e-06, + 8.602978596173e-06,  \
+ 8.621027409390e-06, + 8.637882801850e-06, + 8.653459044581e-06, + 8.667738757140e-06, + 8.680600149091e-06 ]

* Data table for Id-Vd at Vg = 0.34V
.param vd_data_vg0.34=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.34=[ \
+ 9.994420000000e-07, + 1.925400000000e-06, + 2.773000000000e-06, + 3.538300000000e-06, + 4.218600000000e-06,  \
+ 4.814100000000e-06, + 5.327900000000e-06, + 5.766500000000e-06, + 6.137900000000e-06, + 6.450700000000e-06,  \
+ 6.713100000000e-06, + 6.932800000000e-06, + 7.117200000000e-06, + 7.272700000000e-06, + 7.404900000000e-06,  \
+ 7.518600000000e-06, + 7.617400000000e-06, + 7.704600000000e-06, + 7.782300000000e-06, + 7.852400000000e-06,  \
+ 7.916400000000e-06, + 7.975300000000e-06, + 8.030100000000e-06, + 8.081400000000e-06, + 8.129900000000e-06,  \
+ 8.175900000000e-06, + 8.219700000000e-06, + 8.261800000000e-06, + 8.302300000000e-06, + 8.341500000000e-06,  \
+ 8.379400000000e-06, + 8.416300000000e-06, + 8.452200000000e-06, + 8.487300000000e-06, + 8.521700000000e-06,  \
+ 8.555300000000e-06, + 8.588400000000e-06, + 8.620900000000e-06, + 8.652800000000e-06, + 8.684400000000e-06,  \
+ 8.715400000000e-06, + 8.746100000000e-06, + 8.776500000000e-06, + 8.806500000000e-06, + 8.836100000000e-06,  \
+ 8.865500000000e-06, + 8.894600000000e-06, + 8.923500000000e-06, + 8.952100000000e-06, + 8.980500000000e-06,  \
+ 9.008700000000e-06, + 9.036700000000e-06, + 9.064600000000e-06, + 9.092200000000e-06, + 9.119700000000e-06,  \
+ 9.147000000000e-06, + 9.174200000000e-06, + 9.201300000000e-06, + 9.228200000000e-06, + 9.255000000000e-06,  \
+ 9.281600000000e-06, + 9.308200000000e-06, + 9.334600000000e-06, + 9.361000000000e-06, + 9.387300000000e-06,  \
+ 9.413400000000e-06, + 9.439500000000e-06, + 9.465500000000e-06, + 9.491400000000e-06, + 9.517300000000e-06,  \
+ 9.543000000000e-06, + 9.568700000000e-06, + 9.594400000000e-06, + 9.619900000000e-06, + 9.645400000000e-06,  \
+ 9.670900000000e-06, + 9.696300000000e-06, + 9.721600000000e-06, + 9.746900000000e-06, + 9.772200000000e-06 ]

.param id_pred_data_vg0.34=[ \
+ 1.055493412423e-06, + 1.989515876630e-06, + 2.813984756358e-06, + 3.539928875398e-06, + 4.177544178674e-06,  \
+ 4.736216214951e-06, + 5.224554261076e-06, + 5.650414386764e-06, + 6.021007211530e-06, + 6.342821870930e-06,  \
+ 6.621778302360e-06, + 6.863198359497e-06, + 7.071859945427e-06, + 7.252070499817e-06, + 7.407664088532e-06,  \
+ 7.542030652985e-06, + 7.658189097128e-06, + 7.758820647723e-06, + 7.846264161344e-06, + 7.922582881292e-06,  \
+ 7.989558507688e-06, + 8.048741437960e-06, + 8.101478670142e-06, + 8.148931665346e-06, + 8.192099812732e-06,  \
+ 8.231812316808e-06, + 8.268781530205e-06, + 8.303600843647e-06, + 8.336767477886e-06, + 8.368704948225e-06,  \
+ 8.399741655012e-06, + 8.430139860138e-06, + 8.460127883154e-06, + 8.489879983244e-06, + 8.519505809090e-06,  \
+ 8.549126068829e-06, + 8.578788165323e-06, + 8.608576536062e-06, + 8.638497674838e-06, + 8.668592636241e-06,  \
+ 8.698845376784e-06, + 8.729287001188e-06, + 8.759889260546e-06, + 8.790671636234e-06, + 8.821606024867e-06,  \
+ 8.852683567966e-06, + 8.883916580089e-06, + 8.915234939195e-06, + 8.946671659942e-06, + 8.978194273368e-06,  \
+ 9.009788755066e-06, + 9.041415614774e-06, + 9.073076962522e-06, + 9.104750643019e-06, + 9.136398330156e-06,  \
+ 9.167974494630e-06, + 9.199480828102e-06, + 9.230860596290e-06, + 9.262066014344e-06, + 9.293064067606e-06,  \
+ 9.323799386038e-06, + 9.354236080981e-06, + 9.384317154399e-06, + 9.413963416591e-06, + 9.443144472243e-06,  \
+ 9.471763623878e-06, + 9.499792668066e-06, + 9.527135262033e-06, + 9.553748159306e-06, + 9.579518700775e-06,  \
+ 9.604415517970e-06, + 9.628320331103e-06, + 9.651214986661e-06, + 9.672993965069e-06, + 9.693597348814e-06,  \
+ 9.712933679111e-06, + 9.730949095683e-06, + 9.747567200975e-06, + 9.762739746293e-06, + 9.776368824532e-06 ]

* Data table for Id-Vd at Vg = 0.35V
.param vd_data_vg0.35=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.35=[ \
+ 1.067500000000e-06, + 2.063200000000e-06, + 2.981800000000e-06, + 3.818600000000e-06, + 4.570300000000e-06,  \
+ 5.235900000000e-06, + 5.817400000000e-06, + 6.319800000000e-06, + 6.750400000000e-06, + 7.117000000000e-06,  \
+ 7.427800000000e-06, + 7.690300000000e-06, + 7.912000000000e-06, + 8.099600000000e-06, + 8.259300000000e-06,  \
+ 8.396400000000e-06, + 8.515200000000e-06, + 8.619500000000e-06, + 8.711900000000e-06, + 8.794900000000e-06,  \
+ 8.870100000000e-06, + 8.938900000000e-06, + 9.002500000000e-06, + 9.061800000000e-06, + 9.117300000000e-06,  \
+ 9.169800000000e-06, + 9.219700000000e-06, + 9.267300000000e-06, + 9.312900000000e-06, + 9.356800000000e-06,  \
+ 9.399300000000e-06, + 9.440400000000e-06, + 9.480400000000e-06, + 9.519300000000e-06, + 9.557300000000e-06,  \
+ 9.594400000000e-06, + 9.630800000000e-06, + 9.666500000000e-06, + 9.701600000000e-06, + 9.736100000000e-06,  \
+ 9.770100000000e-06, + 9.803600000000e-06, + 9.836700000000e-06, + 9.869400000000e-06, + 9.901600000000e-06,  \
+ 9.933600000000e-06, + 9.965200000000e-06, + 9.996400000000e-06, + 1.002740000000e-05, + 1.005820000000e-05,  \
+ 1.008870000000e-05, + 1.011890000000e-05, + 1.014890000000e-05, + 1.017880000000e-05, + 1.020840000000e-05,  \
+ 1.023780000000e-05, + 1.026710000000e-05, + 1.029610000000e-05, + 1.032510000000e-05, + 1.035380000000e-05,  \
+ 1.038250000000e-05, + 1.041100000000e-05, + 1.043930000000e-05, + 1.046760000000e-05, + 1.049570000000e-05,  \
+ 1.052370000000e-05, + 1.055160000000e-05, + 1.057940000000e-05, + 1.060710000000e-05, + 1.063480000000e-05,  \
+ 1.066230000000e-05, + 1.068970000000e-05, + 1.071710000000e-05, + 1.074440000000e-05, + 1.077160000000e-05,  \
+ 1.079870000000e-05, + 1.082580000000e-05, + 1.085280000000e-05, + 1.087970000000e-05, + 1.090660000000e-05 ]

.param id_pred_data_vg0.35=[ \
+ 1.128153744503e-06, + 2.135361282853e-06, + 3.032336171600e-06, + 3.829123743344e-06, + 4.535140033113e-06,  \
+ 5.159159190953e-06, + 5.709332908737e-06, + 6.193214212544e-06, + 6.617785620620e-06, + 6.989484973019e-06,  \
+ 7.314208924072e-06, + 7.597338699270e-06, + 7.843790008337e-06, + 8.058021412580e-06, + 8.244065065810e-06,  \
+ 8.405562839471e-06, + 8.545771743229e-06, + 8.667600341141e-06, + 8.773649278737e-06, + 8.866240386851e-06,  \
+ 8.947377573350e-06, + 9.018875352922e-06, + 9.082289543585e-06, + 9.138974128291e-06, + 9.190128366754e-06,  \
+ 9.236758560291e-06, + 9.279727455578e-06, + 9.319817181677e-06, + 9.357613125758e-06, + 9.393650179845e-06,  \
+ 9.428352786927e-06, + 9.462112793699e-06, + 9.495192625764e-06, + 9.527830407023e-06, + 9.560229591443e-06,  \
+ 9.592489659553e-06, + 9.624771646486e-06, + 9.657104856160e-06, + 9.689571143099e-06, + 9.722205140861e-06,  \
+ 9.755037463037e-06, + 9.788045572350e-06, + 9.821254134295e-06, + 9.854647214524e-06, + 9.888232671074e-06,  \
+ 9.922007629939e-06, + 9.955892528524e-06, + 9.989923273679e-06, + 1.002405952022e-05, + 1.005830381473e-05,  \
+ 1.009260262435e-05, + 1.012695793179e-05, + 1.016130609059e-05, + 1.019564126182e-05, + 1.022994883897e-05,  \
+ 1.026415920933e-05, + 1.029825398291e-05, + 1.033218850353e-05, + 1.036592153469e-05, + 1.039942399075e-05,  \
+ 1.043260399456e-05, + 1.046543293342e-05, + 1.049786633303e-05, + 1.052981475368e-05, + 1.056122546288e-05,  \
+ 1.059202179022e-05, + 1.062212921170e-05, + 1.065150383511e-05, + 1.068005534762e-05, + 1.070771068044e-05,  \
+ 1.073438196727e-05, + 1.076000167814e-05, + 1.078449696251e-05, + 1.080777112293e-05, + 1.082975859390e-05,  \
+ 1.085037863959e-05, + 1.086955030587e-05, + 1.088721992346e-05, + 1.090331308660e-05, + 1.091770172934e-05 ]

* Data table for Id-Vd at Vg = 0.36V
.param vd_data_vg0.36=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.36=[ \
+ 1.133200000000e-06, + 2.196600000000e-06, + 3.184200000000e-06, + 4.090900000000e-06, + 4.912800000000e-06,  \
+ 5.647900000000e-06, + 6.297300000000e-06, + 6.864700000000e-06, + 7.356300000000e-06, + 7.779500000000e-06,  \
+ 8.141800000000e-06, + 8.450800000000e-06, + 8.713600000000e-06, + 8.937200000000e-06, + 9.128100000000e-06,  \
+ 9.292000000000e-06, + 9.434000000000e-06, + 9.558000000000e-06, + 9.667600000000e-06, + 9.765300000000e-06,  \
+ 9.853400000000e-06, + 9.933700000000e-06, + 1.000730000000e-05, + 1.007560000000e-05, + 1.013930000000e-05,  \
+ 1.019910000000e-05, + 1.025570000000e-05, + 1.030940000000e-05, + 1.036070000000e-05, + 1.040990000000e-05,  \
+ 1.045730000000e-05, + 1.050300000000e-05, + 1.054740000000e-05, + 1.059040000000e-05, + 1.063230000000e-05,  \
+ 1.067320000000e-05, + 1.071310000000e-05, + 1.075220000000e-05, + 1.079060000000e-05, + 1.082830000000e-05,  \
+ 1.086530000000e-05, + 1.090180000000e-05, + 1.093770000000e-05, + 1.097310000000e-05, + 1.100810000000e-05,  \
+ 1.104270000000e-05, + 1.107680000000e-05, + 1.111060000000e-05, + 1.114400000000e-05, + 1.117720000000e-05,  \
+ 1.121000000000e-05, + 1.124250000000e-05, + 1.127480000000e-05, + 1.130680000000e-05, + 1.133860000000e-05,  \
+ 1.137010000000e-05, + 1.140150000000e-05, + 1.143260000000e-05, + 1.146360000000e-05, + 1.149430000000e-05,  \
+ 1.152500000000e-05, + 1.155540000000e-05, + 1.158570000000e-05, + 1.161580000000e-05, + 1.164580000000e-05,  \
+ 1.167570000000e-05, + 1.170540000000e-05, + 1.173500000000e-05, + 1.176450000000e-05, + 1.179390000000e-05,  \
+ 1.182320000000e-05, + 1.185230000000e-05, + 1.188140000000e-05, + 1.191040000000e-05, + 1.193930000000e-05,  \
+ 1.196810000000e-05, + 1.199680000000e-05, + 1.202540000000e-05, + 1.205400000000e-05, + 1.208250000000e-05 ]

.param id_pred_data_vg0.36=[ \
+ 1.197192468680e-06, + 2.274858561577e-06, + 3.242508028052e-06, + 4.109151195735e-06, + 4.883340807282e-06,  \
+ 5.573164526140e-06, + 6.186244136188e-06, + 6.729720043950e-06, + 7.210285330075e-06, + 7.634205394424e-06,  \
+ 8.007257420104e-06, + 8.334842277691e-06, + 8.621909873909e-06, + 8.873025944922e-06, + 9.092390064325e-06,  \
+ 9.283786057495e-06, + 9.450705183554e-06, + 9.596263480489e-06, + 9.723323346407e-06, + 9.834392403718e-06,  \
+ 9.931756248989e-06, + 1.001742268272e-05, + 1.009320865705e-05, + 1.016063906718e-05, + 1.022113792715e-05,  \
+ 1.027589911246e-05, + 1.032596675941e-05, + 1.037223832100e-05, + 1.041545547196e-05, + 1.045629323926e-05,  \
+ 1.049529186275e-05, + 1.053292304277e-05, + 1.056954421074e-05, + 1.060546099325e-05, + 1.064093603418e-05,  \
+ 1.067614990461e-05, + 1.071124101145e-05, + 1.074633266398e-05, + 1.078152483387e-05, + 1.081685695681e-05,  \
+ 1.085236111976e-05, + 1.088805423933e-05, + 1.092396270906e-05, + 1.096006039006e-05, + 1.099637429434e-05,  \
+ 1.103284128476e-05, + 1.106947425797e-05, + 1.110626268201e-05, + 1.114312924983e-05, + 1.118010914070e-05,  \
+ 1.121712055465e-05, + 1.125417737057e-05, + 1.129122811108e-05, + 1.132823545049e-05, + 1.136516184488e-05,  \
+ 1.140198364737e-05, + 1.143863695688e-05, + 1.147511455201e-05, + 1.151132721134e-05, + 1.154725359811e-05,  \
+ 1.158282602773e-05, + 1.161798805697e-05, + 1.165269368357e-05, + 1.168686314486e-05, + 1.172043012048e-05,  \
+ 1.175330457045e-05, + 1.178547699965e-05, + 1.181680680020e-05, + 1.184723934784e-05, + 1.187669258798e-05,  \
+ 1.190509598018e-05, + 1.193236079416e-05, + 1.195840621222e-05, + 1.198312838824e-05, + 1.200645419885e-05,  \
+ 1.202833991556e-05, + 1.204867290653e-05, + 1.206734992593e-05, + 1.208432293424e-05, + 1.209952024510e-05 ]

* Data table for Id-Vd at Vg = 0.37V
.param vd_data_vg0.37=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.37=[ \
+ 1.196600000000e-06, + 2.325300000000e-06, + 3.379800000000e-06, + 4.354500000000e-06, + 5.245000000000e-06,  \
+ 6.048700000000e-06, + 6.765600000000e-06, + 7.398400000000e-06, + 7.952200000000e-06, + 8.433700000000e-06,  \
+ 8.850000000000e-06, + 9.208400000000e-06, + 9.515700000000e-06, + 9.779000000000e-06, + 1.000470000000e-05,  \
+ 1.019890000000e-05, + 1.036700000000e-05, + 1.051380000000e-05, + 1.064290000000e-05, + 1.075770000000e-05,  \
+ 1.086070000000e-05, + 1.095400000000e-05, + 1.103920000000e-05, + 1.111770000000e-05, + 1.119050000000e-05,  \
+ 1.125860000000e-05, + 1.132270000000e-05, + 1.138330000000e-05, + 1.144090000000e-05, + 1.149600000000e-05,  \
+ 1.154880000000e-05, + 1.159950000000e-05, + 1.164860000000e-05, + 1.169610000000e-05, + 1.174220000000e-05,  \
+ 1.178710000000e-05, + 1.183090000000e-05, + 1.187360000000e-05, + 1.191540000000e-05, + 1.195650000000e-05,  \
+ 1.199670000000e-05, + 1.203630000000e-05, + 1.207520000000e-05, + 1.211350000000e-05, + 1.215130000000e-05,  \
+ 1.218850000000e-05, + 1.222530000000e-05, + 1.226170000000e-05, + 1.229760000000e-05, + 1.233320000000e-05,  \
+ 1.236840000000e-05, + 1.240330000000e-05, + 1.243790000000e-05, + 1.247210000000e-05, + 1.250610000000e-05,  \
+ 1.253980000000e-05, + 1.257330000000e-05, + 1.260650000000e-05, + 1.263950000000e-05, + 1.267230000000e-05,  \
+ 1.270490000000e-05, + 1.273730000000e-05, + 1.276950000000e-05, + 1.280160000000e-05, + 1.283350000000e-05,  \
+ 1.286520000000e-05, + 1.289670000000e-05, + 1.292810000000e-05, + 1.295940000000e-05, + 1.299060000000e-05,  \
+ 1.302160000000e-05, + 1.305250000000e-05, + 1.308330000000e-05, + 1.311390000000e-05, + 1.314450000000e-05,  \
+ 1.317500000000e-05, + 1.320530000000e-05, + 1.323560000000e-05, + 1.326570000000e-05, + 1.329580000000e-05 ]

.param id_pred_data_vg0.37=[ \
+ 1.262591831619e-06, + 2.407824067632e-06, + 3.443980385782e-06, + 4.379051970318e-06, + 5.220705497777e-06,  \
+ 5.976271204418e-06, + 6.652783122263e-06, + 7.256902172230e-06, + 7.794950579409e-06, + 8.272930426756e-06,  \
+ 8.696480217623e-06, + 9.070867672563e-06, + 9.401065472048e-06, + 9.691681771073e-06, + 9.946962745744e-06,  \
+ 1.017087721266e-05, + 1.036706460582e-05, + 1.053885105648e-05, + 1.068925204891e-05, + 1.082103044610e-05,  \
+ 1.093669045076e-05, + 1.103845519538e-05, + 1.112836380344e-05, + 1.120815955801e-05, + 1.127946597990e-05,  \
+ 1.134365142207e-05, + 1.140194381151e-05, + 1.145542832091e-05, + 1.150501258962e-05, + 1.155143363576e-05,  \
+ 1.159542469395e-05, + 1.163752167486e-05, + 1.167821723357e-05, + 1.171786738269e-05, + 1.175681718451e-05,  \
+ 1.179530750960e-05, + 1.183351199870e-05, + 1.187162466522e-05, + 1.190975257487e-05, + 1.194796059281e-05,  \
+ 1.198633119202e-05, + 1.202484832902e-05, + 1.206358636409e-05, + 1.210250280565e-05, + 1.214160665768e-05,  \
+ 1.218090630573e-05, + 1.222033755766e-05, + 1.225991029060e-05, + 1.229958565091e-05, + 1.233930925082e-05,  \
+ 1.237908354597e-05, + 1.241886573553e-05, + 1.245861078132e-05, + 1.249826433195e-05, + 1.253780847037e-05,  \
+ 1.257720621652e-05, + 1.261640987650e-05, + 1.265533956030e-05, + 1.269398057048e-05, + 1.273227571801e-05,  \
+ 1.277015808228e-05, + 1.280759392102e-05, + 1.284449210289e-05, + 1.288079423830e-05, + 1.291643402510e-05,  \
+ 1.295131765801e-05, + 1.298540719290e-05, + 1.301861106185e-05, + 1.305083011175e-05, + 1.308199134655e-05,  \
+ 1.311202639044e-05, + 1.314084001933e-05, + 1.316835563557e-05, + 1.319447168498e-05, + 1.321910849583e-05,  \
+ 1.324218152149e-05, + 1.326360590610e-05, + 1.328328009549e-05, + 1.330112561845e-05, + 1.331709063379e-05 ]

* Data table for Id-Vd at Vg = 0.38V
.param vd_data_vg0.38=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.38=[ \
+ 1.257500000000e-06, + 2.449200000000e-06, + 3.568400000000e-06, + 4.609100000000e-06, + 5.566400000000e-06,  \
+ 6.437300000000e-06, + 7.220800000000e-06, + 7.918700000000e-06, + 8.535200000000e-06, + 9.076200000000e-06,  \
+ 9.548400000000e-06, + 9.958400000000e-06, + 1.031310000000e-05, + 1.061910000000e-05, + 1.088290000000e-05,  \
+ 1.111080000000e-05, + 1.130830000000e-05, + 1.148070000000e-05, + 1.163210000000e-05, + 1.176630000000e-05,  \
+ 1.188630000000e-05, + 1.199440000000e-05, + 1.209270000000e-05, + 1.218290000000e-05, + 1.226610000000e-05,  \
+ 1.234360000000e-05, + 1.241610000000e-05, + 1.248430000000e-05, + 1.254900000000e-05, + 1.261050000000e-05,  \
+ 1.266920000000e-05, + 1.272550000000e-05, + 1.277980000000e-05, + 1.283210000000e-05, + 1.288280000000e-05,  \
+ 1.293200000000e-05, + 1.297980000000e-05, + 1.302650000000e-05, + 1.307200000000e-05, + 1.311660000000e-05,  \
+ 1.316020000000e-05, + 1.320300000000e-05, + 1.324510000000e-05, + 1.328640000000e-05, + 1.332710000000e-05,  \
+ 1.336720000000e-05, + 1.340680000000e-05, + 1.344580000000e-05, + 1.348430000000e-05, + 1.352240000000e-05,  \
+ 1.356010000000e-05, + 1.359740000000e-05, + 1.363430000000e-05, + 1.367090000000e-05, + 1.370710000000e-05,  \
+ 1.374300000000e-05, + 1.377870000000e-05, + 1.381400000000e-05, + 1.384910000000e-05, + 1.388390000000e-05,  \
+ 1.391850000000e-05, + 1.395290000000e-05, + 1.398710000000e-05, + 1.402100000000e-05, + 1.405480000000e-05,  \
+ 1.408840000000e-05, + 1.412180000000e-05, + 1.415500000000e-05, + 1.418810000000e-05, + 1.422100000000e-05,  \
+ 1.425380000000e-05, + 1.428640000000e-05, + 1.431890000000e-05, + 1.435120000000e-05, + 1.438340000000e-05,  \
+ 1.441550000000e-05, + 1.444750000000e-05, + 1.447940000000e-05, + 1.451120000000e-05, + 1.454280000000e-05 ]

.param id_pred_data_vg0.38=[ \
+ 1.324447366642e-06, + 2.534262021072e-06, + 3.636576220742e-06, + 4.638337413780e-06, + 5.546330430661e-06,  \
+ 6.367145979311e-06, + 7.107121418812e-06, + 7.772432873026e-06, + 8.368976050406e-06, + 8.902414265322e-06,  \
+ 9.378142058267e-06, + 9.801345295273e-06, + 1.017683767714e-05, + 1.050924052834e-05, + 1.080284673662e-05,  \
+ 1.106171403080e-05, + 1.128956653702e-05, + 1.148991286755e-05, + 1.166595196992e-05, + 1.182064443128e-05,  \
+ 1.195667726279e-05, + 1.207649846037e-05, + 1.218230616360e-05, + 1.227613189258e-05, + 1.235976014868e-05,  \
+ 1.243475169758e-05, + 1.250254990737e-05, + 1.256433679373e-05, + 1.262123623746e-05, + 1.267414372705e-05,  \
+ 1.272390185477e-05, + 1.277115428820e-05, + 1.281649900193e-05, + 1.286041857384e-05, + 1.290331401833e-05,  \
+ 1.294547095313e-05, + 1.298716753809e-05, + 1.302860961005e-05, + 1.306994188781e-05, + 1.311125961365e-05,  \
+ 1.315268924373e-05, + 1.319422444794e-05, + 1.323593347479e-05, + 1.327782221779e-05, + 1.331987223239e-05,  \
+ 1.336206838459e-05, + 1.340442751825e-05, + 1.344688644167e-05, + 1.348939913441e-05, + 1.353197149001e-05,  \
+ 1.357452945740e-05, + 1.361703616567e-05, + 1.365948215607e-05, + 1.370182049868e-05, + 1.374398098051e-05,  \
+ 1.378590619424e-05, + 1.382761103741e-05, + 1.386898213241e-05, + 1.391001593220e-05, + 1.395059516653e-05,  \
+ 1.399072882123e-05, + 1.403033715178e-05, + 1.406932291502e-05, + 1.410767319612e-05, + 1.414527750967e-05,  \
+ 1.418204647052e-05, + 1.421797844159e-05, + 1.425292015483e-05, + 1.428680503523e-05, + 1.431959353795e-05,  \
+ 1.435114183550e-05, + 1.438141538529e-05, + 1.441029193302e-05, + 1.443770161131e-05, + 1.446351416234e-05,  \
+ 1.448770985007e-05, + 1.451015234124e-05, + 1.453073200537e-05, + 1.454943600038e-05, + 1.456612080801e-05 ]

* Data table for Id-Vd at Vg = 0.39V
.param vd_data_vg0.39=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.39=[ \
+ 1.316000000000e-06, + 2.568300000000e-06, + 3.749900000000e-06, + 4.854400000000e-06, + 5.876600000000e-06,  \
+ 6.813000000000e-06, + 7.661900000000e-06, + 8.424300000000e-06, + 9.103500000000e-06, + 9.704600000000e-06,  \
+ 1.023360000000e-05, + 1.069700000000e-05, + 1.110120000000e-05, + 1.145260000000e-05, + 1.175750000000e-05,  \
+ 1.202210000000e-05, + 1.225220000000e-05, + 1.245310000000e-05, + 1.262960000000e-05, + 1.278560000000e-05,  \
+ 1.292480000000e-05, + 1.304970000000e-05, + 1.316290000000e-05, + 1.326620000000e-05, + 1.336120000000e-05,  \
+ 1.344920000000e-05, + 1.353120000000e-05, + 1.360800000000e-05, + 1.368050000000e-05, + 1.374910000000e-05,  \
+ 1.381450000000e-05, + 1.387690000000e-05, + 1.393680000000e-05, + 1.399440000000e-05, + 1.405000000000e-05,  \
+ 1.410390000000e-05, + 1.415610000000e-05, + 1.420690000000e-05, + 1.425650000000e-05, + 1.430480000000e-05,  \
+ 1.435200000000e-05, + 1.439830000000e-05, + 1.444360000000e-05, + 1.448820000000e-05, + 1.453200000000e-05,  \
+ 1.457500000000e-05, + 1.461740000000e-05, + 1.465920000000e-05, + 1.470050000000e-05, + 1.474120000000e-05,  \
+ 1.478140000000e-05, + 1.482120000000e-05, + 1.486050000000e-05, + 1.489940000000e-05, + 1.493800000000e-05,  \
+ 1.497620000000e-05, + 1.501400000000e-05, + 1.505150000000e-05, + 1.508870000000e-05, + 1.512560000000e-05,  \
+ 1.516230000000e-05, + 1.519860000000e-05, + 1.523480000000e-05, + 1.527070000000e-05, + 1.530630000000e-05,  \
+ 1.534180000000e-05, + 1.537700000000e-05, + 1.541210000000e-05, + 1.544700000000e-05, + 1.548160000000e-05,  \
+ 1.551620000000e-05, + 1.555050000000e-05, + 1.558470000000e-05, + 1.561870000000e-05, + 1.565260000000e-05,  \
+ 1.568640000000e-05, + 1.572000000000e-05, + 1.575340000000e-05, + 1.578680000000e-05, + 1.582000000000e-05 ]

.param id_pred_data_vg0.39=[ \
+ 1.382917980663e-06, + 2.654354320839e-06, + 3.820327401627e-06, + 4.886835231446e-06, + 5.859757584403e-06,  \
+ 6.744912680006e-06, + 7.548015273642e-06, + 8.274642750621e-06, + 8.930241383496e-06, + 9.520095773041e-06,  \
+ 1.004934805678e-05, + 1.052291278029e-05, + 1.094553001167e-05, + 1.132172546932e-05, + 1.165576977655e-05,  \
+ 1.195178483613e-05, + 1.221354657901e-05, + 1.244468890945e-05, + 1.264854588953e-05, + 1.282826415263e-05,  \
+ 1.298668743402e-05, + 1.312646621955e-05, + 1.325005130639e-05, + 1.335958979325e-05, + 1.345706550637e-05,  \
+ 1.354430693027e-05, + 1.362286886433e-05, + 1.369416189846e-05, + 1.375945797918e-05, + 1.381979927828e-05,  \
+ 1.387615924614e-05, + 1.392933889292e-05, + 1.398002197675e-05, + 1.402879774105e-05, + 1.407613999618e-05,  \
+ 1.412243946106e-05, + 1.416802140739e-05, + 1.421316301276e-05, + 1.425800943252e-05, + 1.430275588064e-05,  \
+ 1.434748410247e-05, + 1.439227104129e-05, + 1.443716126232e-05, + 1.448220253224e-05, + 1.452736069041e-05,  \
+ 1.457261743781e-05, + 1.461797819502e-05, + 1.466342713684e-05, + 1.470891713325e-05, + 1.475436692999e-05,  \
+ 1.479978094721e-05, + 1.484511893068e-05, + 1.489030026278e-05, + 1.493530005973e-05, + 1.498008377894e-05,  \
+ 1.502457642346e-05, + 1.506873493781e-05, + 1.511249320174e-05, + 1.515584772278e-05, + 1.519868455944e-05,  \
+ 1.524099867311e-05, + 1.528265962406e-05, + 1.532367832624e-05, + 1.536395284347e-05, + 1.540340763313e-05,  \
+ 1.544197464682e-05, + 1.547959307572e-05, + 1.551615445351e-05, + 1.555160464704e-05, + 1.558583844599e-05,  \
+ 1.561883649629e-05, + 1.565041064168e-05, + 1.568051966387e-05, + 1.570907075802e-05, + 1.573600138727e-05,  \
+ 1.576118265803e-05, + 1.578452913236e-05, + 1.580596850545e-05, + 1.582542303368e-05, + 1.584275596542e-05 ]

* Data table for Id-Vd at Vg = 0.40V
.param vd_data_vg0.40=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.40=[ \
+ 1.372100000000e-06, + 2.682600000000e-06, + 3.924200000000e-06, + 5.090300000000e-06, + 6.175300000000e-06,  \
+ 7.175400000000e-06, + 8.088300000000e-06, + 8.914200000000e-06, + 9.655600000000e-06, + 1.031680000000e-05,  \
+ 1.090330000000e-05, + 1.142120000000e-05, + 1.187650000000e-05, + 1.227540000000e-05, + 1.262380000000e-05,  \
+ 1.292790000000e-05, + 1.319330000000e-05, + 1.342570000000e-05, + 1.362990000000e-05, + 1.381050000000e-05,  \
+ 1.397110000000e-05, + 1.411510000000e-05, + 1.424500000000e-05, + 1.436310000000e-05, + 1.447130000000e-05,  \
+ 1.457110000000e-05, + 1.466370000000e-05, + 1.475010000000e-05, + 1.483130000000e-05, + 1.490790000000e-05,  \
+ 1.498050000000e-05, + 1.504970000000e-05, + 1.511580000000e-05, + 1.517920000000e-05, + 1.524020000000e-05,  \
+ 1.529910000000e-05, + 1.535610000000e-05, + 1.541140000000e-05, + 1.546520000000e-05, + 1.551750000000e-05,  \
+ 1.556860000000e-05, + 1.561850000000e-05, + 1.566740000000e-05, + 1.571530000000e-05, + 1.576230000000e-05,  \
+ 1.580850000000e-05, + 1.585390000000e-05, + 1.589860000000e-05, + 1.594270000000e-05, + 1.598610000000e-05,  \
+ 1.602900000000e-05, + 1.607130000000e-05, + 1.611310000000e-05, + 1.615450000000e-05, + 1.619540000000e-05,  \
+ 1.623590000000e-05, + 1.627600000000e-05, + 1.631570000000e-05, + 1.635510000000e-05, + 1.639410000000e-05,  \
+ 1.643280000000e-05, + 1.647120000000e-05, + 1.650940000000e-05, + 1.654720000000e-05, + 1.658480000000e-05,  \
+ 1.662220000000e-05, + 1.665930000000e-05, + 1.669620000000e-05, + 1.673280000000e-05, + 1.676930000000e-05,  \
+ 1.680560000000e-05, + 1.684170000000e-05, + 1.687750000000e-05, + 1.691330000000e-05, + 1.694880000000e-05,  \
+ 1.698420000000e-05, + 1.701940000000e-05, + 1.705450000000e-05, + 1.708950000000e-05, + 1.712430000000e-05 ]

.param id_pred_data_vg0.40=[ \
+ 1.438197796233e-06, + 2.768358681351e-06, + 3.995483421022e-06, + 5.124622839503e-06, + 6.160829070723e-06,  \
+ 7.109163561836e-06, + 7.974672698765e-06, + 8.762364741415e-06, + 9.477190033067e-06, + 1.012405264191e-05,  \
+ 1.070771315426e-05, + 1.123288355302e-05, + 1.170408824692e-05, + 1.212575574755e-05, + 1.250209643331e-05,  \
+ 1.283719786443e-05, + 1.313490189204e-05, + 1.339890834060e-05, + 1.363266324915e-05, + 1.383943745168e-05,  \
+ 1.402221962053e-05, + 1.418387968442e-05, + 1.432698045392e-05, + 1.445389701985e-05, + 1.456685731682e-05,  \
+ 1.466779584007e-05, + 1.475849036069e-05, + 1.484050924773e-05, + 1.491529634222e-05, + 1.498409255873e-05,  \
+ 1.504796997324e-05, + 1.510787289590e-05, + 1.516460950370e-05, + 1.521888225398e-05, + 1.527128933958e-05,  \
+ 1.532223555841e-05, + 1.537217274745e-05, + 1.542138779769e-05, + 1.547013434902e-05, + 1.551863970235e-05,  \
+ 1.556697789056e-05, + 1.561528893944e-05, + 1.566360606375e-05, + 1.571197892190e-05, + 1.576043032401e-05,  \
+ 1.580894044309e-05, + 1.585749978403e-05, + 1.590607396793e-05, + 1.595461275429e-05, + 1.600310315553e-05,  \
+ 1.605147237569e-05, + 1.609966158867e-05, + 1.614766002604e-05, + 1.619537906663e-05, + 1.624281039767e-05,  \
+ 1.628987272852e-05, + 1.633650417716e-05, + 1.638266236114e-05, + 1.642828208787e-05, + 1.647333192523e-05,  \
+ 1.651774540733e-05, + 1.656144417211e-05, + 1.660438974795e-05, + 1.664649113081e-05, + 1.668768054515e-05,  \
+ 1.672791477176e-05, + 1.676711532127e-05, + 1.680514622421e-05, + 1.684203220066e-05, + 1.687759249762e-05,  \
+ 1.691180934358e-05, + 1.694455946563e-05, + 1.697578158200e-05, + 1.700536206044e-05, + 1.703321549940e-05,  \
+ 1.705926828436e-05, + 1.708344621875e-05, + 1.710557167826e-05, + 1.712566234346e-05, + 1.714355312288e-05 ]

* Data table for Id-Vd at Vg = 0.41V
.param vd_data_vg0.41=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.41=[ \
+ 1.425800000000e-06, + 2.792100000000e-06, + 4.091400000000e-06, + 5.316800000000e-06, + 6.462600000000e-06,  \
+ 7.524400000000e-06, + 8.499600000000e-06, + 9.387800000000e-06, + 1.019060000000e-05, + 1.091160000000e-05,  \
+ 1.155580000000e-05, + 1.212880000000e-05, + 1.263630000000e-05, + 1.308410000000e-05, + 1.347810000000e-05,  \
+ 1.382390000000e-05, + 1.412730000000e-05, + 1.439380000000e-05, + 1.462850000000e-05, + 1.483600000000e-05,  \
+ 1.502060000000e-05, + 1.518570000000e-05, + 1.533430000000e-05, + 1.546900000000e-05, + 1.559200000000e-05,  \
+ 1.570500000000e-05, + 1.580950000000e-05, + 1.590660000000e-05, + 1.599740000000e-05, + 1.608290000000e-05,  \
+ 1.616360000000e-05, + 1.624010000000e-05, + 1.631310000000e-05, + 1.638280000000e-05, + 1.644970000000e-05,  \
+ 1.651410000000e-05, + 1.657630000000e-05, + 1.663640000000e-05, + 1.669480000000e-05, + 1.675140000000e-05,  \
+ 1.680660000000e-05, + 1.686050000000e-05, + 1.691310000000e-05, + 1.696450000000e-05, + 1.701490000000e-05,  \
+ 1.706440000000e-05, + 1.711300000000e-05, + 1.716070000000e-05, + 1.720770000000e-05, + 1.725400000000e-05,  \
+ 1.729960000000e-05, + 1.734460000000e-05, + 1.738900000000e-05, + 1.743280000000e-05, + 1.747620000000e-05,  \
+ 1.751910000000e-05, + 1.756150000000e-05, + 1.760350000000e-05, + 1.764510000000e-05, + 1.768630000000e-05,  \
+ 1.772710000000e-05, + 1.776760000000e-05, + 1.780780000000e-05, + 1.784760000000e-05, + 1.788720000000e-05,  \
+ 1.792650000000e-05, + 1.796550000000e-05, + 1.800420000000e-05, + 1.804270000000e-05, + 1.808100000000e-05,  \
+ 1.811900000000e-05, + 1.815680000000e-05, + 1.819440000000e-05, + 1.823190000000e-05, + 1.826910000000e-05,  \
+ 1.830610000000e-05, + 1.834300000000e-05, + 1.837970000000e-05, + 1.841620000000e-05, + 1.845260000000e-05 ]

.param id_pred_data_vg0.41=[ \
+ 1.490507129347e-06, + 2.876606886275e-06, + 4.162367113167e-06, + 5.351967993192e-06, + 6.449643842643e-06,  \
+ 7.459767221007e-06, + 8.386695408262e-06, + 9.234870085493e-06, + 1.000876181934e-05, + 1.071283040801e-05,  \
+ 1.135148137109e-05, + 1.192910625832e-05, + 1.245005310921e-05, + 1.291857595788e-05, + 1.333876862191e-05,  \
+ 1.371465972625e-05, + 1.405013324984e-05, + 1.434887919459e-05, + 1.461441941501e-05, + 1.485015527578e-05,  \
+ 1.505920488853e-05, + 1.524453458842e-05, + 1.540892750199e-05, + 1.555493508931e-05, + 1.568493462401e-05,  \
+ 1.580104712048e-05, + 1.590523981577e-05, + 1.599927578354e-05, + 1.608470323845e-05, + 1.616300723981e-05,  \
+ 1.623533269594e-05, + 1.630287035368e-05, + 1.636643428355e-05, + 1.642690447625e-05, + 1.648494981055e-05,  \
+ 1.654114370467e-05, + 1.659592395299e-05, + 1.664970761340e-05, + 1.670278237725e-05, + 1.675536041148e-05,  \
+ 1.680764751654e-05, + 1.685977607849e-05, + 1.691178254987e-05, + 1.696380029898e-05, + 1.701577093627e-05,  \
+ 1.706773815386e-05, + 1.711965807772e-05, + 1.717155799270e-05, + 1.722333345242e-05, + 1.727497146931e-05,  \
+ 1.732639117108e-05, + 1.737759856042e-05, + 1.742847547575e-05, + 1.747902824718e-05, + 1.752914849931e-05,  \
+ 1.757879828801e-05, + 1.762792544469e-05, + 1.767648598616e-05, + 1.772440635250e-05, + 1.777162106009e-05,  \
+ 1.781807301086e-05, + 1.786372926290e-05, + 1.790851549231e-05, + 1.795238233171e-05, + 1.799522315196e-05,  \
+ 1.803701077733e-05, + 1.807760683732e-05, + 1.811705551518e-05, + 1.815517585783e-05, + 1.819192966650e-05,  \
+ 1.822722944780e-05, + 1.826102903578e-05, + 1.829317763622e-05, + 1.832360208937e-05, + 1.835228476921e-05,  \
+ 1.837905809225e-05, + 1.840387825723e-05, + 1.842660742113e-05, + 1.844717646236e-05, + 1.846553059295e-05 ]

* Data table for Id-Vd at Vg = 0.42V
.param vd_data_vg0.42=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.42=[ \
+ 1.477200000000e-06, + 2.896900000000e-06, + 4.251600000000e-06, + 5.534000000000e-06, + 6.738400000000e-06,  \
+ 7.859900000000e-06, + 8.895700000000e-06, + 9.844600000000e-06, + 1.070780000000e-05, + 1.148810000000e-05,  \
+ 1.218970000000e-05, + 1.281800000000e-05, + 1.337830000000e-05, + 1.387620000000e-05, + 1.431720000000e-05,  \
+ 1.470670000000e-05, + 1.505020000000e-05, + 1.535320000000e-05, + 1.562080000000e-05, + 1.585780000000e-05,  \
+ 1.606860000000e-05, + 1.625710000000e-05, + 1.642650000000e-05, + 1.657970000000e-05, + 1.671920000000e-05,  \
+ 1.684690000000e-05, + 1.696450000000e-05, + 1.707360000000e-05, + 1.717520000000e-05, + 1.727040000000e-05,  \
+ 1.736000000000e-05, + 1.744470000000e-05, + 1.752520000000e-05, + 1.760190000000e-05, + 1.767520000000e-05,  \
+ 1.774560000000e-05, + 1.781340000000e-05, + 1.787880000000e-05, + 1.794200000000e-05, + 1.800340000000e-05,  \
+ 1.806300000000e-05, + 1.812100000000e-05, + 1.817750000000e-05, + 1.823280000000e-05, + 1.828680000000e-05,  \
+ 1.833970000000e-05, + 1.839160000000e-05, + 1.844260000000e-05, + 1.849260000000e-05, + 1.854190000000e-05,  \
+ 1.859040000000e-05, + 1.863810000000e-05, + 1.868520000000e-05, + 1.873170000000e-05, + 1.877760000000e-05,  \
+ 1.882290000000e-05, + 1.886770000000e-05, + 1.891200000000e-05, + 1.895590000000e-05, + 1.899930000000e-05,  \
+ 1.904230000000e-05, + 1.908500000000e-05, + 1.912720000000e-05, + 1.916910000000e-05, + 1.921070000000e-05,  \
+ 1.925190000000e-05, + 1.929280000000e-05, + 1.933340000000e-05, + 1.937380000000e-05, + 1.941390000000e-05,  \
+ 1.945370000000e-05, + 1.949330000000e-05, + 1.953260000000e-05, + 1.957180000000e-05, + 1.961070000000e-05,  \
+ 1.964930000000e-05, + 1.968780000000e-05, + 1.972610000000e-05, + 1.976430000000e-05, + 1.980220000000e-05 ]

.param id_pred_data_vg0.42=[ \
+ 1.540072262287e-06, + 2.979459532071e-06, + 4.321387968957e-06, + 5.569222266786e-06, + 6.726470019203e-06,  \
+ 7.796786958352e-06, + 8.783935190877e-06, + 9.691776940599e-06, + 1.052426261595e-05, + 1.128541116486e-05,  \
+ 1.197927929752e-05, + 1.260994904442e-05, + 1.318145434198e-05, + 1.369787787553e-05, + 1.416324666934e-05,  \
+ 1.458141021430e-05, + 1.495618918852e-05, + 1.529136919999e-05, + 1.559047443152e-05, + 1.585691788932e-05,  \
+ 1.609399449080e-05, + 1.630475890124e-05, + 1.649215642828e-05, + 1.665891031735e-05, + 1.680747845967e-05,  \
+ 1.694025268080e-05, + 1.705934046186e-05, + 1.716661616229e-05, + 1.726395552396e-05, + 1.735279984132e-05,  \
+ 1.743463853927e-05, + 1.751062110998e-05, + 1.758186230290e-05, + 1.764929715137e-05, + 1.771365423338e-05,  \
+ 1.777566445526e-05, + 1.783584259101e-05, + 1.789465117326e-05, + 1.795246465917e-05, + 1.800957834348e-05,  \
+ 1.806619362469e-05, + 1.812246722693e-05, + 1.817849009967e-05, + 1.823440281441e-05, + 1.829019674915e-05,  \
+ 1.834582930314e-05, + 1.840139073465e-05, + 1.845677266829e-05, + 1.851199798693e-05, + 1.856693415903e-05,  \
+ 1.862166707724e-05, + 1.867595317890e-05, + 1.872986405942e-05, + 1.878331459011e-05, + 1.883624081529e-05,  \
+ 1.888854778372e-05, + 1.894023353088e-05, + 1.899119466543e-05, + 1.904142482090e-05, + 1.909080165206e-05,  \
+ 1.913929740113e-05, + 1.918689282320e-05, + 1.923345422256e-05, + 1.927902339958e-05, + 1.932337163453e-05,  \
+ 1.936663589731e-05, + 1.940857655427e-05, + 1.944926130818e-05, + 1.948852917849e-05, + 1.952632628672e-05,  \
+ 1.956255387995e-05, + 1.959720393643e-05, + 1.963015036381e-05, + 1.966129930224e-05, + 1.969059258045e-05,  \
+ 1.971790748939e-05, + 1.974321728994e-05, + 1.976639417990e-05, + 1.978730693736e-05, + 1.980595698114e-05 ]

* Data table for Id-Vd at Vg = 0.43V
.param vd_data_vg0.43=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.43=[ \
+ 1.526300000000e-06, + 2.997200000000e-06, + 4.404900000000e-06, + 5.742200000000e-06, + 7.002900000000e-06,  \
+ 8.182100000000e-06, + 9.276500000000e-06, + 1.028470000000e-05, + 1.120700000000e-05, + 1.204560000000e-05,  \
+ 1.280430000000e-05, + 1.348770000000e-05, + 1.410110000000e-05, + 1.464960000000e-05, + 1.513860000000e-05,  \
+ 1.557320000000e-05, + 1.595870000000e-05, + 1.630030000000e-05, + 1.660310000000e-05, + 1.687190000000e-05,  \
+ 1.711120000000e-05, + 1.732530000000e-05, + 1.751750000000e-05, + 1.769110000000e-05, + 1.784880000000e-05,  \
+ 1.799280000000e-05, + 1.812510000000e-05, + 1.824740000000e-05, + 1.836090000000e-05, + 1.846690000000e-05,  \
+ 1.856630000000e-05, + 1.866010000000e-05, + 1.874880000000e-05, + 1.883310000000e-05, + 1.891350000000e-05,  \
+ 1.899040000000e-05, + 1.906430000000e-05, + 1.913530000000e-05, + 1.920390000000e-05, + 1.927030000000e-05,  \
+ 1.933460000000e-05, + 1.939710000000e-05, + 1.945790000000e-05, + 1.951720000000e-05, + 1.957510000000e-05,  \
+ 1.963170000000e-05, + 1.968710000000e-05, + 1.974140000000e-05, + 1.979470000000e-05, + 1.984700000000e-05,  \
+ 1.989850000000e-05, + 1.994920000000e-05, + 1.999910000000e-05, + 2.004830000000e-05, + 2.009680000000e-05,  \
+ 2.014470000000e-05, + 2.019200000000e-05, + 2.023870000000e-05, + 2.028490000000e-05, + 2.033060000000e-05,  \
+ 2.037590000000e-05, + 2.042070000000e-05, + 2.046500000000e-05, + 2.050900000000e-05, + 2.055260000000e-05,  \
+ 2.059580000000e-05, + 2.063870000000e-05, + 2.068120000000e-05, + 2.072350000000e-05, + 2.076540000000e-05,  \
+ 2.080700000000e-05, + 2.084840000000e-05, + 2.088950000000e-05, + 2.093040000000e-05, + 2.097100000000e-05,  \
+ 2.101130000000e-05, + 2.105150000000e-05, + 2.109140000000e-05, + 2.113110000000e-05, + 2.117060000000e-05 ]

.param id_pred_data_vg0.43=[ \
+ 1.587107253727e-06, + 3.077284782194e-06, + 4.472975560930e-06, + 5.776832695119e-06, + 6.991661211941e-06,  \
+ 8.120491693262e-06, + 9.166457748506e-06, + 1.013291068375e-05, + 1.102326481487e-05, + 1.184113934869e-05,  \
+ 1.259019372810e-05, + 1.327412581304e-05, + 1.389674922393e-05, + 1.446189722628e-05, + 1.497341436334e-05,  \
+ 1.543503371067e-05, + 1.585054640600e-05, + 1.622359923203e-05, + 1.655781183217e-05, + 1.685663009994e-05,  \
+ 1.712339348160e-05, + 1.736125836032e-05, + 1.757326339430e-05, + 1.776232849807e-05, + 1.793104456738e-05,  \
+ 1.808190048905e-05, + 1.821724734327e-05, + 1.833911490394e-05, + 1.844945349148e-05, + 1.855002265074e-05,  \
+ 1.864236095571e-05, + 1.872773165815e-05, + 1.880751166027e-05, + 1.888261795102e-05, + 1.895403984236e-05,  \
+ 1.902249612613e-05, + 1.908866179292e-05, + 1.915302505950e-05, + 1.921607825352e-05, + 1.927813136717e-05,  \
+ 1.933945259225e-05, + 1.940024689247e-05, + 1.946066575329e-05, + 1.952078353497e-05, + 1.958064312930e-05,  \
+ 1.964029368537e-05, + 1.969968157937e-05, + 1.975885767024e-05, + 1.981769713893e-05, + 1.987622272281e-05,  \
+ 1.993432222662e-05, + 1.999195781536e-05, + 2.004903577472e-05, + 2.010554082517e-05, + 2.016136713792e-05,  \
+ 2.021646563662e-05, + 2.027076068771e-05, + 2.032425531070e-05, + 2.037678863417e-05, + 2.042836131295e-05,  \
+ 2.047894420684e-05, + 2.052842442936e-05, + 2.057677076664e-05, + 2.062392653897e-05, + 2.066985234705e-05,  \
+ 2.071443108434e-05, + 2.075762724417e-05, + 2.079941594275e-05, + 2.083969993691e-05, + 2.087842549372e-05,  \
+ 2.091546572046e-05, + 2.095083415043e-05, + 2.098439459587e-05, + 2.101606984070e-05, + 2.104583472828e-05,  \
+ 2.107354237523e-05, + 2.109918450515e-05, + 2.112256253895e-05, + 2.114372151482e-05, + 2.116245741490e-05 ]

* Data table for Id-Vd at Vg = 0.44V
.param vd_data_vg0.44=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.44=[ \
+ 1.573200000000e-06, + 3.093000000000e-06, + 4.551600000000e-06, + 5.941400000000e-06, + 7.256300000000e-06,  \
+ 8.491100000000e-06, + 9.642300000000e-06, + 1.070800000000e-05, + 1.168790000000e-05, + 1.258380000000e-05,  \
+ 1.339880000000e-05, + 1.413710000000e-05, + 1.480350000000e-05, + 1.540300000000e-05, + 1.594060000000e-05,  \
+ 1.642140000000e-05, + 1.685020000000e-05, + 1.723200000000e-05, + 1.757190000000e-05, + 1.787460000000e-05,  \
+ 1.814470000000e-05, + 1.838640000000e-05, + 1.860350000000e-05, + 1.879950000000e-05, + 1.897720000000e-05,  \
+ 1.913910000000e-05, + 1.928760000000e-05, + 1.942440000000e-05, + 1.955110000000e-05, + 1.966900000000e-05,  \
+ 1.977930000000e-05, + 1.988290000000e-05, + 1.998070000000e-05, + 2.007340000000e-05, + 2.016150000000e-05,  \
+ 2.024550000000e-05, + 2.032600000000e-05, + 2.040320000000e-05, + 2.047760000000e-05, + 2.054940000000e-05,  \
+ 2.061880000000e-05, + 2.068610000000e-05, + 2.075140000000e-05, + 2.081500000000e-05, + 2.087700000000e-05,  \
+ 2.093750000000e-05, + 2.099660000000e-05, + 2.105450000000e-05, + 2.111120000000e-05, + 2.116680000000e-05,  \
+ 2.122150000000e-05, + 2.127520000000e-05, + 2.132800000000e-05, + 2.138000000000e-05, + 2.143130000000e-05,  \
+ 2.148180000000e-05, + 2.153170000000e-05, + 2.158090000000e-05, + 2.162950000000e-05, + 2.167760000000e-05,  \
+ 2.172520000000e-05, + 2.177220000000e-05, + 2.181880000000e-05, + 2.186490000000e-05, + 2.191050000000e-05,  \
+ 2.195580000000e-05, + 2.200070000000e-05, + 2.204520000000e-05, + 2.208930000000e-05, + 2.213310000000e-05,  \
+ 2.217660000000e-05, + 2.221980000000e-05, + 2.226270000000e-05, + 2.230530000000e-05, + 2.234760000000e-05,  \
+ 2.238960000000e-05, + 2.243140000000e-05, + 2.247300000000e-05, + 2.251430000000e-05, + 2.255540000000e-05 ]

.param id_pred_data_vg0.44=[ \
+ 1.631817576708e-06, + 3.170417621732e-06, + 4.617573868018e-06, + 5.975256790407e-06, + 7.245667802636e-06,  \
+ 8.431213209406e-06, + 9.534508571960e-06, + 1.055830740370e-05, + 1.150565381977e-05, + 1.237961987499e-05,  \
+ 1.318349233770e-05, + 1.392070669681e-05, + 1.459472892748e-05, + 1.520913458080e-05, + 1.576754839334e-05,  \
+ 1.627361285500e-05, + 1.673096361628e-05, + 1.714321842883e-05, + 1.751393770974e-05, + 1.784656342352e-05,  \
+ 1.814450792153e-05, + 1.841101882746e-05, + 1.864921439847e-05, + 1.886208134238e-05, + 1.905237877509e-05,  \
+ 1.922278592247e-05, + 1.937568857102e-05, + 1.951347367140e-05, + 1.963806796994e-05, + 1.975142440642e-05,  \
+ 1.985525195778e-05, + 1.995104830712e-05, + 2.004018653679e-05, + 2.012384262343e-05, + 2.020300235017e-05,  \
+ 2.027856098721e-05, + 2.035126948613e-05, + 2.042176027317e-05, + 2.049055285170e-05, + 2.055801451206e-05,  \
+ 2.062448900688e-05, + 2.069019210467e-05, + 2.075534041069e-05, + 2.081999395159e-05, + 2.088427463605e-05,  \
+ 2.094819770718e-05, + 2.101176065480e-05, + 2.107497886755e-05, + 2.113771777658e-05, + 2.119999953720e-05,  \
+ 2.126172385033e-05, + 2.132285240805e-05, + 2.138336258213e-05, + 2.144307647541e-05, + 2.150198033632e-05,  \
+ 2.156000322429e-05, + 2.161706208426e-05, + 2.167313694372e-05, + 2.172810025513e-05, + 2.178195136366e-05,  \
+ 2.183461561799e-05, + 2.188603357354e-05, + 2.193617663579e-05, + 2.198494039476e-05, + 2.203229705628e-05,  \
+ 2.207819576142e-05, + 2.212258958025e-05, + 2.216543274699e-05, + 2.220660466264e-05, + 2.224610980193e-05,  \
+ 2.228385597846e-05, + 2.231979276985e-05, + 2.235381762148e-05, + 2.238589462650e-05, + 2.241593347208e-05,  \
+ 2.244383933430e-05, + 2.246960473713e-05, + 2.249310771731e-05, + 2.251424313727e-05, + 2.253299171571e-05 ]

* Data table for Id-Vd at Vg = 0.45V
.param vd_data_vg0.45=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.45=[ \
+ 1.618000000000e-06, + 3.184600000000e-06, + 4.691700000000e-06, + 6.132000000000e-06, + 7.498900000000e-06,  \
+ 8.787300000000e-06, + 9.993300000000e-06, + 1.111460000000e-05, + 1.215080000000e-05, + 1.310270000000e-05,  \
+ 1.397310000000e-05, + 1.476560000000e-05, + 1.548470000000e-05, + 1.613520000000e-05, + 1.672180000000e-05,  \
+ 1.724930000000e-05, + 1.772240000000e-05, + 1.814580000000e-05, + 1.852440000000e-05, + 1.886280000000e-05,  \
+ 1.916560000000e-05, + 1.943700000000e-05, + 1.968100000000e-05, + 1.990120000000e-05, + 2.010070000000e-05,  \
+ 2.028240000000e-05, + 2.044860000000e-05, + 2.060130000000e-05, + 2.074250000000e-05, + 2.087350000000e-05,  \
+ 2.099570000000e-05, + 2.111020000000e-05, + 2.121790000000e-05, + 2.131970000000e-05, + 2.141620000000e-05,  \
+ 2.150800000000e-05, + 2.159570000000e-05, + 2.167970000000e-05, + 2.176030000000e-05, + 2.183790000000e-05,  \
+ 2.191280000000e-05, + 2.198530000000e-05, + 2.205550000000e-05, + 2.212370000000e-05, + 2.219000000000e-05,  \
+ 2.225470000000e-05, + 2.231780000000e-05, + 2.237940000000e-05, + 2.243970000000e-05, + 2.249880000000e-05,  \
+ 2.255680000000e-05, + 2.261370000000e-05, + 2.266960000000e-05, + 2.272450000000e-05, + 2.277860000000e-05,  \
+ 2.283190000000e-05, + 2.288450000000e-05, + 2.293630000000e-05, + 2.298750000000e-05, + 2.303800000000e-05,  \
+ 2.308790000000e-05, + 2.313720000000e-05, + 2.318600000000e-05, + 2.323430000000e-05, + 2.328220000000e-05,  \
+ 2.332950000000e-05, + 2.337640000000e-05, + 2.342290000000e-05, + 2.346910000000e-05, + 2.351480000000e-05,  \
+ 2.356010000000e-05, + 2.360510000000e-05, + 2.364980000000e-05, + 2.369420000000e-05, + 2.373820000000e-05,  \
+ 2.378200000000e-05, + 2.382550000000e-05, + 2.386870000000e-05, + 2.391160000000e-05, + 2.395430000000e-05 ]

.param id_pred_data_vg0.45=[ \
+ 1.674392406130e-06, + 3.259199729655e-06, + 4.755594563903e-06, + 6.164967198856e-06, + 7.488935079891e-06,  \
+ 8.729373221286e-06, + 9.888352506096e-06, + 1.096818596125e-05, + 1.197134843096e-05, + 1.290061627515e-05,  \
+ 1.375882697175e-05, + 1.454907964217e-05, + 1.527450433059e-05, + 1.593844397576e-05, + 1.654430634517e-05,  \
+ 1.709552132525e-05, + 1.759562626830e-05, + 1.804814441130e-05, + 1.845657105150e-05, + 1.882430806290e-05,  \
+ 1.915480905154e-05, + 1.945140233147e-05, + 1.971717290871e-05, + 1.995530154090e-05, + 2.016862708842e-05,  \
+ 2.035992758465e-05, + 2.053179989161e-05, + 2.068666100968e-05, + 2.082672886900e-05, + 2.095400050166e-05,  \
+ 2.107037820679e-05, + 2.117754891515e-05, + 2.127693602233e-05, + 2.136987022823e-05, + 2.145757498511e-05,  \
+ 2.154092668206e-05, + 2.162084165320e-05, + 2.169804771256e-05, + 2.177304941142e-05, + 2.184640034102e-05,  \
+ 2.191844054323e-05, + 2.198950365710e-05, + 2.205973112723e-05, + 2.212931285612e-05, + 2.219833604613e-05,  \
+ 2.226685377536e-05, + 2.233486655314e-05, + 2.240238420200e-05, + 2.246931111586e-05, + 2.253564525745e-05,  \
+ 2.260127999762e-05, + 2.266619470902e-05, + 2.273028007039e-05, + 2.279345018906e-05, + 2.285562732141e-05,  \
+ 2.291673619766e-05, + 2.297674887814e-05, + 2.303551642399e-05, + 2.309305444214e-05, + 2.314927114639e-05,  \
+ 2.320411465917e-05, + 2.325755944184e-05, + 2.330946470465e-05, + 2.335990080610e-05, + 2.340867922612e-05,  \
+ 2.345590102777e-05, + 2.350140635826e-05, + 2.354521391680e-05, + 2.358724021178e-05, + 2.362744126003e-05,  \
+ 2.366574997723e-05, + 2.370212838287e-05, + 2.373647279455e-05, + 2.376878823270e-05, + 2.379900342930e-05,  \
+ 2.382697217399e-05, + 2.385268799117e-05, + 2.387608736171e-05, + 2.389706549366e-05, + 2.391557354713e-05 ]

* Data table for Id-Vd at Vg = 0.46V
.param vd_data_vg0.46=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.46=[ \
+ 1.660700000000e-06, + 3.272000000000e-06, + 4.825600000000e-06, + 6.314200000000e-06, + 7.731000000000e-06,  \
+ 9.070900000000e-06, + 1.032970000000e-05, + 1.150500000000e-05, + 1.259560000000e-05, + 1.360230000000e-05,  \
+ 1.452710000000e-05, + 1.537310000000e-05, + 1.614440000000e-05, + 1.684560000000e-05, + 1.748120000000e-05,  \
+ 1.805570000000e-05, + 1.857370000000e-05, + 1.903980000000e-05, + 1.945830000000e-05, + 1.983400000000e-05,  \
+ 2.017110000000e-05, + 2.047410000000e-05, + 2.074680000000e-05, + 2.099310000000e-05, + 2.121620000000e-05,  \
+ 2.141920000000e-05, + 2.160470000000e-05, + 2.177490000000e-05, + 2.193190000000e-05, + 2.207730000000e-05,  \
+ 2.221250000000e-05, + 2.233890000000e-05, + 2.245750000000e-05, + 2.256920000000e-05, + 2.267490000000e-05,  \
+ 2.277520000000e-05, + 2.287070000000e-05, + 2.296190000000e-05, + 2.304930000000e-05, + 2.313320000000e-05,  \
+ 2.321410000000e-05, + 2.329210000000e-05, + 2.336750000000e-05, + 2.344070000000e-05, + 2.351170000000e-05,  \
+ 2.358080000000e-05, + 2.364810000000e-05, + 2.371370000000e-05, + 2.377790000000e-05, + 2.384060000000e-05,  \
+ 2.390210000000e-05, + 2.396230000000e-05, + 2.402140000000e-05, + 2.407950000000e-05, + 2.413660000000e-05,  \
+ 2.419280000000e-05, + 2.424810000000e-05, + 2.430260000000e-05, + 2.435640000000e-05, + 2.440950000000e-05,  \
+ 2.446180000000e-05, + 2.451360000000e-05, + 2.456470000000e-05, + 2.461530000000e-05, + 2.466530000000e-05,  \
+ 2.471480000000e-05, + 2.476380000000e-05, + 2.481240000000e-05, + 2.486050000000e-05, + 2.490820000000e-05,  \
+ 2.495540000000e-05, + 2.500230000000e-05, + 2.504880000000e-05, + 2.509500000000e-05, + 2.514080000000e-05,  \
+ 2.518630000000e-05, + 2.523150000000e-05, + 2.527640000000e-05, + 2.532100000000e-05, + 2.536530000000e-05 ]

.param id_pred_data_vg0.46=[ \
+ 1.714990648907e-06, + 3.343930875417e-06, + 4.887438408332e-06, + 6.346412701532e-06, + 7.721937436145e-06,  \
+ 9.015401301440e-06, + 1.022838987410e-05, + 1.136274659075e-05, + 1.242053069291e-05, + 1.340410963167e-05,  \
+ 1.431595112081e-05, + 1.515874697361e-05, + 1.593537643203e-05, + 1.664890762186e-05, + 1.730248986860e-05,  \
+ 1.789942034520e-05, + 1.844299564254e-05, + 1.893665496027e-05, + 1.938377645274e-05, + 1.978781365324e-05,  \
+ 2.015209662204e-05, + 2.048002381343e-05, + 2.077474418911e-05, + 2.103944483679e-05, + 2.127713923983e-05,  \
+ 2.149067324353e-05, + 2.168277795136e-05, + 2.185596938943e-05, + 2.201260242146e-05, + 2.215495915152e-05,  \
+ 2.228493380244e-05, + 2.240441506729e-05, + 2.251494726806e-05, + 2.261805624585e-05, + 2.271493358421e-05,  \
+ 2.280684420839e-05, + 2.289455696882e-05, + 2.297902712598e-05, + 2.306080976268e-05, + 2.314057492185e-05,  \
+ 2.321865369595e-05, + 2.329544346139e-05, + 2.337117854040e-05, + 2.344603824895e-05, + 2.352017691010e-05,  \
+ 2.359362952120e-05, + 2.366643791902e-05, + 2.373857132625e-05, + 2.381001180765e-05, + 2.388069151493e-05,  \
+ 2.395049519691e-05, + 2.401942139841e-05, + 2.408737807855e-05, + 2.415420633042e-05, + 2.421986500849e-05,  \
+ 2.428429521387e-05, + 2.434737831209e-05, + 2.440911703161e-05, + 2.446933951433e-05, + 2.452806365909e-05,  \
+ 2.458521328663e-05, + 2.464073520969e-05, + 2.469454931997e-05, + 2.474665874615e-05, + 2.479701015545e-05,  \
+ 2.484546756023e-05, + 2.489212762157e-05, + 2.493688429240e-05, + 2.497970384866e-05, + 2.502051502233e-05,  \
+ 2.505931122869e-05, + 2.509606245439e-05, + 2.513065381208e-05, + 2.516306674806e-05, + 2.519325062167e-05,  \
+ 2.522112714360e-05, + 2.524666248064e-05, + 2.526976626541e-05, + 2.529044981202e-05, + 2.530856290832e-05 ]

* Data table for Id-Vd at Vg = 0.47V
.param vd_data_vg0.47=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.47=[ \
+ 1.701500000000e-06, + 3.355400000000e-06, + 4.953500000000e-06, + 6.488200000000e-06, + 7.953000000000e-06,  \
+ 9.342300000000e-06, + 1.065200000000e-05, + 1.187930000000e-05, + 1.302290000000e-05, + 1.408280000000e-05,  \
+ 1.506070000000e-05, + 1.595930000000e-05, + 1.678230000000e-05, + 1.753370000000e-05, + 1.821810000000e-05,  \
+ 1.883970000000e-05, + 1.940300000000e-05, + 1.991230000000e-05, + 2.037180000000e-05, + 2.078590000000e-05,  \
+ 2.115880000000e-05, + 2.149490000000e-05, + 2.179810000000e-05, + 2.207220000000e-05, + 2.232070000000e-05,  \
+ 2.254670000000e-05, + 2.275310000000e-05, + 2.294220000000e-05, + 2.311630000000e-05, + 2.327730000000e-05,  \
+ 2.342680000000e-05, + 2.356610000000e-05, + 2.369660000000e-05, + 2.381920000000e-05, + 2.393480000000e-05,  \
+ 2.404430000000e-05, + 2.414830000000e-05, + 2.424740000000e-05, + 2.434210000000e-05, + 2.443290000000e-05,  \
+ 2.452010000000e-05, + 2.460410000000e-05, + 2.468520000000e-05, + 2.476360000000e-05, + 2.483970000000e-05,  \
+ 2.491350000000e-05, + 2.498520000000e-05, + 2.505520000000e-05, + 2.512340000000e-05, + 2.519000000000e-05,  \
+ 2.525510000000e-05, + 2.531890000000e-05, + 2.538140000000e-05, + 2.544270000000e-05, + 2.550300000000e-05,  \
+ 2.556220000000e-05, + 2.562040000000e-05, + 2.567780000000e-05, + 2.573430000000e-05, + 2.578990000000e-05,  \
+ 2.584490000000e-05, + 2.589910000000e-05, + 2.595260000000e-05, + 2.600550000000e-05, + 2.605780000000e-05,  \
+ 2.610950000000e-05, + 2.616070000000e-05, + 2.621140000000e-05, + 2.626150000000e-05, + 2.631120000000e-05,  \
+ 2.636050000000e-05, + 2.640930000000e-05, + 2.645770000000e-05, + 2.650570000000e-05, + 2.655330000000e-05,  \
+ 2.660060000000e-05, + 2.664750000000e-05, + 2.669410000000e-05, + 2.674030000000e-05, + 2.678630000000e-05 ]

.param id_pred_data_vg0.47=[ \
+ 1.753766118782e-06, + 3.424868918955e-06, + 5.013476475142e-06, + 6.520015886053e-06, + 7.945130346343e-06,  \
+ 9.289737499785e-06, + 1.055498636561e-05, + 1.174232689664e-05, + 1.285341670155e-05, + 1.389013923472e-05,  \
+ 1.485472152126e-05, + 1.574943889864e-05, + 1.657694985624e-05, + 1.733990007779e-05, + 1.804132953112e-05,  \
+ 1.868421211839e-05, + 1.927175318997e-05, + 1.980723085580e-05, + 2.029392402619e-05, + 2.073519572150e-05,  \
+ 2.113436748914e-05, + 2.149475432816e-05, + 2.181963558542e-05, + 2.211217302829e-05, + 2.237549233541e-05,  \
+ 2.261246714625e-05, + 2.282602566993e-05, + 2.301877480932e-05, + 2.319320512470e-05, + 2.335163517273e-05,  \
+ 2.349627073272e-05, + 2.362900413573e-05, + 2.375158030191e-05, + 2.386567823123e-05, + 2.397263087914e-05,  \
+ 2.407364838291e-05, + 2.416987408651e-05, + 2.426217281027e-05, + 2.435130983940e-05, + 2.443791599944e-05,  \
+ 2.452247645124e-05, + 2.460545372742e-05, + 2.468707334629e-05, + 2.476763620507e-05, + 2.484725646354e-05,  \
+ 2.492599465768e-05, + 2.500391681679e-05, + 2.508098899852e-05, + 2.515723506804e-05, + 2.523251532693e-05,  \
+ 2.530687583203e-05, + 2.538009212003e-05, + 2.545214232669e-05, + 2.552297373768e-05, + 2.559235435911e-05,  \
+ 2.566036186181e-05, + 2.572682282334e-05, + 2.579164305644e-05, + 2.585480691778e-05, + 2.591621378087e-05,  \
+ 2.597582770250e-05, + 2.603357148473e-05, + 2.608940900245e-05, + 2.614331431687e-05, + 2.619523493195e-05,  \
+ 2.624507294968e-05, + 2.629288141179e-05, + 2.633860087371e-05, + 2.638221583766e-05, + 2.642362742336e-05,  \
+ 2.646288405231e-05, + 2.649984788150e-05, + 2.653457868291e-05, + 2.656700453372e-05, + 2.659707206476e-05,  \
+ 2.662472412339e-05, + 2.664995110536e-05, + 2.667268730875e-05, + 2.669283694559e-05, + 2.671040128917e-05 ]

* Data table for Id-Vd at Vg = 0.48V
.param vd_data_vg0.48=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.48=[ \
+ 1.740400000000e-06, + 3.435000000000e-06, + 5.075600000000e-06, + 6.654500000000e-06, + 8.165200000000e-06,  \
+ 9.602000000000e-06, + 1.096060000000e-05, + 1.223810000000e-05, + 1.343280000000e-05, + 1.454450000000e-05,  \
+ 1.557430000000e-05, + 1.652440000000e-05, + 1.739820000000e-05, + 1.819940000000e-05, + 1.893220000000e-05,  \
+ 1.960080000000e-05, + 2.020940000000e-05, + 2.076220000000e-05, + 2.126330000000e-05, + 2.171670000000e-05,  \
+ 2.212670000000e-05, + 2.249720000000e-05, + 2.283240000000e-05, + 2.313590000000e-05, + 2.341130000000e-05,  \
+ 2.366190000000e-05, + 2.389070000000e-05, + 2.410030000000e-05, + 2.429300000000e-05, + 2.447090000000e-05,  \
+ 2.463580000000e-05, + 2.478920000000e-05, + 2.493250000000e-05, + 2.506690000000e-05, + 2.519340000000e-05,  \
+ 2.531290000000e-05, + 2.542610000000e-05, + 2.553370000000e-05, + 2.563640000000e-05, + 2.573450000000e-05,  \
+ 2.582860000000e-05, + 2.591900000000e-05, + 2.600620000000e-05, + 2.609030000000e-05, + 2.617160000000e-05,  \
+ 2.625050000000e-05, + 2.632710000000e-05, + 2.640150000000e-05, + 2.647400000000e-05, + 2.654470000000e-05,  \
+ 2.661380000000e-05, + 2.668130000000e-05, + 2.674740000000e-05, + 2.681220000000e-05, + 2.687570000000e-05,  \
+ 2.693810000000e-05, + 2.699940000000e-05, + 2.705960000000e-05, + 2.711900000000e-05, + 2.717740000000e-05,  \
+ 2.723500000000e-05, + 2.729180000000e-05, + 2.734780000000e-05, + 2.740310000000e-05, + 2.745780000000e-05,  \
+ 2.751180000000e-05, + 2.756520000000e-05, + 2.761800000000e-05, + 2.767030000000e-05, + 2.772200000000e-05,  \
+ 2.777330000000e-05, + 2.782400000000e-05, + 2.787440000000e-05, + 2.792420000000e-05, + 2.797370000000e-05,  \
+ 2.802280000000e-05, + 2.807140000000e-05, + 2.811980000000e-05, + 2.816770000000e-05, + 2.821530000000e-05 ]

.param id_pred_data_vg0.48=[ \
+ 1.790846145013e-06, + 3.502264444251e-06, + 5.134036618983e-06, + 6.686164997518e-06, + 8.158932178048e-06,  \
+ 9.552805277053e-06, + 1.086859221687e-05, + 1.210729475133e-05, + 1.327022124315e-05, + 1.435891317669e-05,  \
+ 1.537515738164e-05, + 1.632103929296e-05, + 1.719879423035e-05, + 1.801089674700e-05, + 1.876003298094e-05,  \
+ 1.944901072420e-05, + 2.008087103604e-05, + 2.065864100587e-05, + 2.118558018992e-05, + 2.166484919144e-05,  \
+ 2.209982325439e-05, + 2.249372104416e-05, + 2.284984395374e-05, + 2.317139238585e-05, + 2.346145993215e-05,  \
+ 2.372312243097e-05, + 2.395930154307e-05, + 2.417272829916e-05, + 2.436600916553e-05, + 2.454164714436e-05,  \
+ 2.470194398484e-05, + 2.484885742888e-05, + 2.498440764612e-05, + 2.511024751584e-05, + 2.522799804865e-05,  \
+ 2.533892024076e-05, + 2.544425435190e-05, + 2.554497841629e-05, + 2.564198301116e-05, + 2.573597594164e-05,  \
+ 2.582751483715e-05, + 2.591708514956e-05, + 2.600506435556e-05, + 2.609166884213e-05, + 2.617711907078e-05,  \
+ 2.626149922435e-05, + 2.634485132148e-05, + 2.642726583872e-05, + 2.650859220012e-05, + 2.658885387063e-05,  \
+ 2.666797281563e-05, + 2.674581759493e-05, + 2.682233232917e-05, + 2.689738910703e-05, + 2.697083837120e-05,  \
+ 2.704263810301e-05, + 2.711273089517e-05, + 2.718096548051e-05, + 2.724724370637e-05, + 2.731159547693e-05,  \
+ 2.737381862971e-05, + 2.743401571934e-05, + 2.749201768893e-05, + 2.754785120487e-05, + 2.760145234788e-05,  \
+ 2.765275312413e-05, + 2.770183233224e-05, + 2.774854539894e-05, + 2.779295879009e-05, + 2.783501877275e-05,  \
+ 2.787464487483e-05, + 2.791190257994e-05, + 2.794672567688e-05, + 2.797911285597e-05, + 2.800893707899e-05,  \
+ 2.803626455716e-05, + 2.806106360367e-05, + 2.808323588397e-05, + 2.810273672367e-05, + 2.811962040141e-05 ]

* Data table for Id-Vd at Vg = 0.49V
.param vd_data_vg0.49=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.49=[ \
+ 1.777500000000e-06, + 3.510900000000e-06, + 5.192100000000e-06, + 6.813300000000e-06, + 8.367900000000e-06,  \
+ 9.850200000000e-06, + 1.125590000000e-05, + 1.258180000000e-05, + 1.382590000000e-05, + 1.498780000000e-05,  \
+ 1.606810000000e-05, + 1.706860000000e-05, + 1.799220000000e-05, + 1.884250000000e-05, + 1.962320000000e-05,  \
+ 2.033850000000e-05, + 2.099230000000e-05, + 2.158880000000e-05, + 2.213170000000e-05, + 2.262520000000e-05,  \
+ 2.307300000000e-05, + 2.347910000000e-05, + 2.384750000000e-05, + 2.418180000000e-05, + 2.448570000000e-05,  \
+ 2.476240000000e-05, + 2.501510000000e-05, + 2.524650000000e-05, + 2.545920000000e-05, + 2.565530000000e-05,  \
+ 2.583690000000e-05, + 2.600550000000e-05, + 2.616270000000e-05, + 2.630990000000e-05, + 2.644810000000e-05,  \
+ 2.657840000000e-05, + 2.670160000000e-05, + 2.681840000000e-05, + 2.692960000000e-05, + 2.703570000000e-05,  \
+ 2.713720000000e-05, + 2.723460000000e-05, + 2.732820000000e-05, + 2.741840000000e-05, + 2.750550000000e-05,  \
+ 2.758970000000e-05, + 2.767140000000e-05, + 2.775070000000e-05, + 2.782780000000e-05, + 2.790280000000e-05,  \
+ 2.797600000000e-05, + 2.804750000000e-05, + 2.811740000000e-05, + 2.818580000000e-05, + 2.825280000000e-05,  \
+ 2.831850000000e-05, + 2.838290000000e-05, + 2.844630000000e-05, + 2.850860000000e-05, + 2.856990000000e-05,  \
+ 2.863020000000e-05, + 2.868970000000e-05, + 2.874830000000e-05, + 2.880610000000e-05, + 2.886320000000e-05,  \
+ 2.891960000000e-05, + 2.897530000000e-05, + 2.903030000000e-05, + 2.908480000000e-05, + 2.913870000000e-05,  \
+ 2.919200000000e-05, + 2.924480000000e-05, + 2.929700000000e-05, + 2.934880000000e-05, + 2.940020000000e-05,  \
+ 2.945110000000e-05, + 2.950160000000e-05, + 2.955170000000e-05, + 2.960130000000e-05, + 2.965070000000e-05 ]

.param id_pred_data_vg0.49=[ \
+ 1.826332882047e-06, + 3.576319722924e-06, + 5.249405221548e-06, + 6.845245370641e-06, + 8.363750384888e-06,  \
+ 9.805042936932e-06, + 1.116956089390e-05, + 1.245797728188e-05, + 1.367123899399e-05, + 1.481056096964e-05,  \
+ 1.587741397088e-05, + 1.687349402346e-05, + 1.780082820915e-05, + 1.866151054855e-05, + 1.945812764461e-05,  \
+ 2.019316656515e-05, + 2.086943510221e-05, + 2.148984553060e-05, + 2.205749937275e-05, + 2.257547312183e-05,  \
+ 2.304701083631e-05, + 2.347531364649e-05, + 2.386360712990e-05, + 2.421518904157e-05, + 2.453312845319e-05,  \
+ 2.482056384906e-05, + 2.508041317924e-05, + 2.531562960939e-05, + 2.552888130595e-05, + 2.572273588157e-05,  \
+ 2.589958974568e-05, + 2.606167690828e-05, + 2.621104264108e-05, + 2.634954260429e-05, + 2.647880937729e-05,  \
+ 2.660033118445e-05, + 2.671539332368e-05, + 2.682516293135e-05, + 2.693057336728e-05, + 2.703243517317e-05,  \
+ 2.713143454457e-05, + 2.722804274526e-05, + 2.732271277637e-05, + 2.741577191046e-05, + 2.750741878117e-05,  \
+ 2.759777191386e-05, + 2.768695194391e-05, + 2.777494140901e-05, + 2.786174263747e-05, + 2.794732790790e-05,  \
+ 2.803153187415e-05, + 2.811432204908e-05, + 2.819558420015e-05, + 2.827518539561e-05, + 2.835296400008e-05,  \
+ 2.842893183697e-05, + 2.850291897630e-05, + 2.857478648366e-05, + 2.864454640076e-05, + 2.871203250834e-05,  \
+ 2.877717328374e-05, + 2.883998829930e-05, + 2.890041119826e-05, + 2.895830431953e-05, + 2.901373754867e-05,  \
+ 2.906671928940e-05, + 2.911711329944e-05, + 2.916499113780e-05, + 2.921024835814e-05, + 2.925294975284e-05,  \
+ 2.929305683210e-05, + 2.933056064649e-05, + 2.936549870356e-05, + 2.939768222859e-05, + 2.942730407085e-05,  \
+ 2.945424988866e-05, + 2.947844528535e-05, + 2.950002155558e-05, + 2.951881560875e-05, + 2.953480579890e-05 ]

* Data table for Id-Vd at Vg = 0.50V
.param vd_data_vg0.50=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.50=[ \
+ 1.812900000000e-06, + 3.583400000000e-06, + 5.303300000000e-06, + 6.964900000000e-06, + 8.561500000000e-06,  \
+ 1.008760000000e-05, + 1.153840000000e-05, + 1.291080000000e-05, + 1.420270000000e-05, + 1.541310000000e-05,  \
+ 1.654250000000e-05, + 1.759220000000e-05, + 1.856470000000e-05, + 1.946310000000e-05, + 2.029110000000e-05,  \
+ 2.105260000000e-05, + 2.175140000000e-05, + 2.239140000000e-05, + 2.297640000000e-05, + 2.351020000000e-05,  \
+ 2.399650000000e-05, + 2.443900000000e-05, + 2.484170000000e-05, + 2.520800000000e-05, + 2.554160000000e-05,  \
+ 2.584580000000e-05, + 2.612380000000e-05, + 2.637850000000e-05, + 2.661250000000e-05, + 2.682810000000e-05,  \
+ 2.702750000000e-05, + 2.721250000000e-05, + 2.738480000000e-05, + 2.754570000000e-05, + 2.769660000000e-05,  \
+ 2.783850000000e-05, + 2.797240000000e-05, + 2.809930000000e-05, + 2.821970000000e-05, + 2.833430000000e-05,  \
+ 2.844380000000e-05, + 2.854860000000e-05, + 2.864920000000e-05, + 2.874590000000e-05, + 2.883910000000e-05,  \
+ 2.892910000000e-05, + 2.901620000000e-05, + 2.910060000000e-05, + 2.918260000000e-05, + 2.926230000000e-05,  \
+ 2.933990000000e-05, + 2.941550000000e-05, + 2.948940000000e-05, + 2.956160000000e-05, + 2.963220000000e-05,  \
+ 2.970140000000e-05, + 2.976930000000e-05, + 2.983580000000e-05, + 2.990120000000e-05, + 2.996550000000e-05,  \
+ 3.002870000000e-05, + 3.009100000000e-05, + 3.015230000000e-05, + 3.021270000000e-05, + 3.027230000000e-05,  \
+ 3.033120000000e-05, + 3.038920000000e-05, + 3.044660000000e-05, + 3.050330000000e-05, + 3.055930000000e-05,  \
+ 3.061480000000e-05, + 3.066960000000e-05, + 3.072400000000e-05, + 3.077770000000e-05, + 3.083100000000e-05,  \
+ 3.088380000000e-05, + 3.093610000000e-05, + 3.098800000000e-05, + 3.103940000000e-05, + 3.109050000000e-05 ]

.param id_pred_data_vg0.50=[ \
+ 1.860323245637e-06, + 3.647225094028e-06, + 5.359851638786e-06, + 6.997558521107e-06, + 8.559935668018e-06,  \
+ 1.004681456834e-05, + 1.145832429756e-05, + 1.279478077777e-05, + 1.405684059137e-05, + 1.524537074147e-05,  \
+ 1.636155851884e-05, + 1.740682579111e-05, + 1.838286829297e-05, + 1.929158868734e-05, + 2.013519770117e-05,  \
+ 2.091606846079e-05, + 2.163675890188e-05, + 2.229998266557e-05, + 2.290866963449e-05, + 2.346580149606e-05,  \
+ 2.397453979938e-05, + 2.443799545290e-05, + 2.485939388862e-05, + 2.524186740629e-05, + 2.558860796853e-05,  \
+ 2.590280695586e-05, + 2.618744321808e-05, + 2.644544758368e-05, + 2.667966509762e-05, + 2.689269458642e-05,  \
+ 2.708714644541e-05, + 2.726527396590e-05, + 2.742935554124e-05, + 2.758126283879e-05, + 2.772278567136e-05,  \
+ 2.785562071949e-05, + 2.798110232106e-05, + 2.810044257785e-05, + 2.821484486049e-05, + 2.832504687831e-05,  \
+ 2.843195346941e-05, + 2.853596888599e-05, + 2.863778005121e-05, + 2.873764518881e-05, + 2.883585875679e-05,  \
+ 2.893256358220e-05, + 2.902785396145e-05, + 2.912182593718e-05, + 2.921445277025e-05, + 2.930564733106e-05,  \
+ 2.939528945717e-05, + 2.948334484245e-05, + 2.956969216029e-05, + 2.965416235384e-05, + 2.973667033075e-05,  \
+ 2.981702855323e-05, + 2.989525328303e-05, + 2.997108887939e-05, + 3.004454498296e-05, + 3.011544467881e-05,  \
+ 3.018382562004e-05, + 3.024951111001e-05, + 3.031254054804e-05, + 3.037279704586e-05, + 3.043032884307e-05,  \
+ 3.048505539482e-05, + 3.053697666473e-05, + 3.058610745938e-05, + 3.063234496949e-05, + 3.067577781621e-05,  \
+ 3.071645907767e-05, + 3.075426095165e-05, + 3.078922200075e-05, + 3.082140698098e-05, + 3.085072967224e-05,  \
+ 3.087723962381e-05, + 3.090086640441e-05, + 3.092168510193e-05, + 3.093961360719e-05, + 3.095472056884e-05 ]

* Data table for Id-Vd at Vg = 0.51V
.param vd_data_vg0.51=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.51=[ \
+ 1.846600000000e-06, + 3.652500000000e-06, + 5.409400000000e-06, + 7.109600000000e-06, + 8.746500000000e-06,  \
+ 1.031440000000e-05, + 1.180860000000e-05, + 1.322580000000e-05, + 1.456360000000e-05, + 1.582100000000e-05,  \
+ 1.699790000000e-05, + 1.809550000000e-05, + 1.911570000000e-05, + 2.006150000000e-05, + 2.093610000000e-05,  \
+ 2.174320000000e-05, + 2.248650000000e-05, + 2.316980000000e-05, + 2.379680000000e-05, + 2.437100000000e-05,  \
+ 2.489610000000e-05, + 2.537580000000e-05, + 2.581340000000e-05, + 2.621280000000e-05, + 2.657720000000e-05,  \
+ 2.691020000000e-05, + 2.721480000000e-05, + 2.749400000000e-05, + 2.775060000000e-05, + 2.798700000000e-05,  \
+ 2.820540000000e-05, + 2.840790000000e-05, + 2.859630000000e-05, + 2.877200000000e-05, + 2.893650000000e-05,  \
+ 2.909090000000e-05, + 2.923640000000e-05, + 2.937390000000e-05, + 2.950430000000e-05, + 2.962810000000e-05,  \
+ 2.974620000000e-05, + 2.985890000000e-05, + 2.996700000000e-05, + 3.007070000000e-05, + 3.017040000000e-05,  \
+ 3.026660000000e-05, + 3.035950000000e-05, + 3.044940000000e-05, + 3.053650000000e-05, + 3.062110000000e-05,  \
+ 3.070340000000e-05, + 3.078350000000e-05, + 3.086160000000e-05, + 3.093780000000e-05, + 3.101230000000e-05,  \
+ 3.108510000000e-05, + 3.115650000000e-05, + 3.122650000000e-05, + 3.129510000000e-05, + 3.136250000000e-05,  \
+ 3.142870000000e-05, + 3.149390000000e-05, + 3.155800000000e-05, + 3.162110000000e-05, + 3.168340000000e-05,  \
+ 3.174470000000e-05, + 3.180530000000e-05, + 3.186500000000e-05, + 3.192400000000e-05, + 3.198230000000e-05,  \
+ 3.204000000000e-05, + 3.209700000000e-05, + 3.215340000000e-05, + 3.220920000000e-05, + 3.226440000000e-05,  \
+ 3.231910000000e-05, + 3.237330000000e-05, + 3.242710000000e-05, + 3.248030000000e-05, + 3.253310000000e-05 ]

.param id_pred_data_vg0.51=[ \
+ 1.892898144433e-06, + 3.715129569173e-06, + 5.465596768772e-06, + 7.143389084376e-06, + 8.747848914936e-06,  \
+ 1.027851743856e-05, + 1.173523080070e-05, + 1.311803935096e-05, + 1.442729058908e-05, + 1.566361024743e-05,  \
+ 1.682783913566e-05, + 1.792117254809e-05, + 1.894498069305e-05, + 1.990093151107e-05, + 2.079102487187e-05,  \
+ 2.161731943488e-05, + 2.238222645246e-05, + 2.308830851689e-05, + 2.373817857006e-05, + 2.433483023196e-05,  \
+ 2.488124278898e-05, + 2.538046988775e-05, + 2.583563116787e-05, + 2.624984190334e-05, + 2.662631959538e-05,  \
+ 2.696820025449e-05, + 2.727853716351e-05, + 2.756032423349e-05, + 2.781645518553e-05, + 2.804968753480e-05,  \
+ 2.826263822499e-05, + 2.845774870366e-05, + 2.863728142984e-05, + 2.880337473471e-05, + 2.895796351368e-05,  \
+ 2.910271170549e-05, + 2.923921958427e-05, + 2.936879624031e-05, + 2.949263805931e-05, + 2.961173013318e-05,  \
+ 2.972692076582e-05, + 2.983885889989e-05, + 2.994820439199e-05, + 3.005522215972e-05, + 3.016035334440e-05,  \
+ 3.026371879969e-05, + 3.036551068362e-05, + 3.046575933695e-05, + 3.056443907553e-05, + 3.066157296416e-05,  \
+ 3.075703396462e-05, + 3.085066884523e-05, + 3.094240801147e-05, + 3.103207061940e-05, + 3.111963033007e-05,  \
+ 3.120479726931e-05, + 3.128752745397e-05, + 3.136764236842e-05, + 3.144518319459e-05, + 3.151986747980e-05,  \
+ 3.159167852573e-05, + 3.166057897033e-05, + 3.172648739564e-05, + 3.178937360644e-05, + 3.184916186001e-05,  \
+ 3.190589341102e-05, + 3.195953340764e-05, + 3.201009836630e-05, + 3.205757180694e-05, + 3.210192408005e-05,  \
+ 3.214314685465e-05, + 3.218138474040e-05, + 3.221652521461e-05, + 3.224863416108e-05, + 3.227768047509e-05,  \
+ 3.230375179555e-05, + 3.232683669921e-05, + 3.234689000237e-05, + 3.236391788960e-05, + 3.237798810005e-05 ]

* Data table for Id-Vd at Vg = 0.52V
.param vd_data_vg0.52=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.52=[ \
+ 1.878800000000e-06, + 3.718400000000e-06, + 5.510600000000e-06, + 7.247800000000e-06, + 8.923200000000e-06,  \
+ 1.053120000000e-05, + 1.206700000000e-05, + 1.352720000000e-05, + 1.490930000000e-05, + 1.621200000000e-05,  \
+ 1.743500000000e-05, + 1.857900000000e-05, + 1.964590000000e-05, + 2.063790000000e-05, + 2.155830000000e-05,  \
+ 2.241030000000e-05, + 2.319760000000e-05, + 2.392390000000e-05, + 2.459260000000e-05, + 2.520720000000e-05,  \
+ 2.577130000000e-05, + 2.628830000000e-05, + 2.676160000000e-05, + 2.719470000000e-05, + 2.759100000000e-05,  \
+ 2.795370000000e-05, + 2.828600000000e-05, + 2.859100000000e-05, + 2.887140000000e-05, + 2.912970000000e-05,  \
+ 2.936840000000e-05, + 2.958960000000e-05, + 2.979510000000e-05, + 2.998660000000e-05, + 3.016560000000e-05,  \
+ 3.033350000000e-05, + 3.049140000000e-05, + 3.064040000000e-05, + 3.078130000000e-05, + 3.091510000000e-05,  \
+ 3.104230000000e-05, + 3.116360000000e-05, + 3.127960000000e-05, + 3.139080000000e-05, + 3.149750000000e-05,  \
+ 3.160030000000e-05, + 3.169940000000e-05, + 3.179510000000e-05, + 3.188770000000e-05, + 3.197750000000e-05,  \
+ 3.206470000000e-05, + 3.214950000000e-05, + 3.223200000000e-05, + 3.231250000000e-05, + 3.239100000000e-05,  \
+ 3.246780000000e-05, + 3.254290000000e-05, + 3.261640000000e-05, + 3.268840000000e-05, + 3.275910000000e-05,  \
+ 3.282850000000e-05, + 3.289670000000e-05, + 3.296370000000e-05, + 3.302970000000e-05, + 3.309460000000e-05,  \
+ 3.315860000000e-05, + 3.322170000000e-05, + 3.328390000000e-05, + 3.334530000000e-05, + 3.340600000000e-05,  \
+ 3.346590000000e-05, + 3.352510000000e-05, + 3.358360000000e-05, + 3.364150000000e-05, + 3.369880000000e-05,  \
+ 3.375550000000e-05, + 3.381160000000e-05, + 3.386720000000e-05, + 3.392230000000e-05, + 3.397690000000e-05 ]

.param id_pred_data_vg0.52=[ \
+ 1.924123062054e-06, + 3.780175466090e-06, + 5.566840991378e-06, + 7.283008890226e-06, + 8.927780436352e-06,  \
+ 1.050046237651e-05, + 1.200064201839e-05, + 1.342811272480e-05, + 1.478297926951e-05, + 1.606558362255e-05,  \
+ 1.727650393150e-05, + 1.841661287472e-05, + 1.948718811036e-05, + 2.048954309430e-05, + 2.142538432963e-05,  \
+ 2.229661447927e-05, + 2.310542462510e-05, + 2.385415253229e-05, + 2.454537228914e-05, + 2.518175751902e-05,  \
+ 2.576617553132e-05, + 2.630161165143e-05, + 2.679114753846e-05, + 2.723776444327e-05, + 2.764477721939e-05,  \
+ 2.801517170155e-05, + 2.835207233147e-05, + 2.865855843993e-05, + 2.893750446674e-05, + 2.919180042227e-05,  \
+ 2.942410952528e-05, + 2.963701495901e-05, + 2.983289225085e-05, + 3.001399076311e-05, + 3.018232855538e-05,  \
+ 3.033970511751e-05, + 3.048786064028e-05, + 3.062817238970e-05, + 3.076204608078e-05, + 3.089044475928e-05,  \
+ 3.101442722254e-05, + 3.113468672382e-05, + 3.125188020931e-05, + 3.136642830214e-05, + 3.147881689074e-05,  \
+ 3.158920429996e-05, + 3.169774718117e-05, + 3.180461120792e-05, + 3.190972820448e-05, + 3.201308936696e-05,  \
+ 3.211459646991e-05, + 3.221414313884e-05, + 3.231163394958e-05, + 3.240690246457e-05, + 3.249973506172e-05,  \
+ 3.259007848101e-05, + 3.267766576755e-05, + 3.276246563473e-05, + 3.284432965302e-05, + 3.292312248959e-05,  \
+ 3.299873031210e-05, + 3.307120248792e-05, + 3.314026922453e-05, + 3.320605261251e-05, + 3.326850564918e-05,  \
+ 3.332747815875e-05, + 3.338309437822e-05, + 3.343530639540e-05, + 3.348412654304e-05, + 3.352952444402e-05,  \
+ 3.357158846484e-05, + 3.361030801898e-05, + 3.364578835317e-05, + 3.367794233782e-05, + 3.370683043613e-05,  \
+ 3.373254221515e-05, + 3.375500877155e-05, + 3.377427136002e-05, + 3.379043802852e-05, + 3.380342095625e-05 ]

* Data table for Id-Vd at Vg = 0.53V
.param vd_data_vg0.53=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.53=[ \
+ 1.909500000000e-06, + 3.781300000000e-06, + 5.607300000000e-06, + 7.379700000000e-06, + 9.092000000000e-06,  \
+ 1.073830000000e-05, + 1.231410000000e-05, + 1.381560000000e-05, + 1.524030000000e-05, + 1.658660000000e-05,  \
+ 1.785420000000e-05, + 1.904340000000e-05, + 2.015550000000e-05, + 2.119280000000e-05, + 2.215800000000e-05,  \
+ 2.305420000000e-05, + 2.388490000000e-05, + 2.465360000000e-05, + 2.536360000000e-05, + 2.601850000000e-05,  \
+ 2.662160000000e-05, + 2.717610000000e-05, + 2.768540000000e-05, + 2.815280000000e-05, + 2.858160000000e-05,  \
+ 2.897490000000e-05, + 2.933590000000e-05, + 2.966770000000e-05, + 2.997300000000e-05, + 3.025440000000e-05,  \
+ 3.051450000000e-05, + 3.075540000000e-05, + 3.097910000000e-05, + 3.118740000000e-05, + 3.138200000000e-05,  \
+ 3.156420000000e-05, + 3.173530000000e-05, + 3.189660000000e-05, + 3.204890000000e-05, + 3.219310000000e-05,  \
+ 3.233020000000e-05, + 3.246060000000e-05, + 3.258510000000e-05, + 3.270430000000e-05, + 3.281850000000e-05,  \
+ 3.292820000000e-05, + 3.303390000000e-05, + 3.313580000000e-05, + 3.323430000000e-05, + 3.332970000000e-05,  \
+ 3.342210000000e-05, + 3.351180000000e-05, + 3.359910000000e-05, + 3.368400000000e-05, + 3.376680000000e-05,  \
+ 3.384770000000e-05, + 3.392660000000e-05, + 3.400390000000e-05, + 3.407950000000e-05, + 3.415360000000e-05,  \
+ 3.422630000000e-05, + 3.429760000000e-05, + 3.436770000000e-05, + 3.443660000000e-05, + 3.450440000000e-05,  \
+ 3.457120000000e-05, + 3.463690000000e-05, + 3.470170000000e-05, + 3.476560000000e-05, + 3.482860000000e-05,  \
+ 3.489090000000e-05, + 3.495230000000e-05, + 3.501310000000e-05, + 3.507310000000e-05, + 3.513250000000e-05,  \
+ 3.519120000000e-05, + 3.524930000000e-05, + 3.530690000000e-05, + 3.536390000000e-05, + 3.542030000000e-05 ]

.param id_pred_data_vg0.53=[ \
+ 1.954048930202e-06, + 3.842466685455e-06, + 5.663767224178e-06, + 7.416644948535e-06, + 9.100011084229e-06,  \
+ 1.071297941962e-05, + 1.225489817443e-05, + 1.372536877170e-05, + 1.512419868959e-05, + 1.645154115977e-05,  \
+ 1.770773858880e-05, + 1.889345236123e-05, + 2.000963810133e-05, + 2.105737454258e-05, + 2.203820622526e-05,  \
+ 2.295378362760e-05, + 2.380606398219e-05, + 2.459718991304e-05, + 2.532957340009e-05, + 2.600572770461e-05,  \
+ 2.662843500730e-05, + 2.720046031754e-05, + 2.772483014269e-05, + 2.820451743901e-05, + 2.864266207325e-05,  \
+ 2.904229302658e-05, + 2.940654587292e-05, + 2.973854891025e-05, + 3.004118399986e-05, + 3.031734813703e-05,  \
+ 3.056989575271e-05, + 3.080143127590e-05, + 3.101446643996e-05, + 3.121125060716e-05, + 3.139402688248e-05,  \
+ 3.156473336276e-05, + 3.172510332661e-05, + 3.187676004018e-05, + 3.202113082807e-05, + 3.215938631911e-05,  \
+ 3.229255467886e-05, + 3.242148435675e-05, + 3.254690527683e-05, + 3.266934276326e-05, + 3.278927833890e-05,  \
+ 3.290698849014e-05, + 3.302267577965e-05, + 3.313637687825e-05, + 3.324820776470e-05, + 3.335806832183e-05,  \
+ 3.346601028170e-05, + 3.357179841259e-05, + 3.367532037373e-05, + 3.377644781722e-05, + 3.387491560716e-05,  \
+ 3.397073305678e-05, + 3.406362360693e-05, + 3.415338956984e-05, + 3.423996888159e-05, + 3.432325611357e-05,  \
+ 3.440309468715e-05, + 3.447937648161e-05, + 3.455200894678e-05, + 3.462099004537e-05, + 3.468630529824e-05,  \
+ 3.474792240013e-05, + 3.480580955511e-05, + 3.485988112516e-05, + 3.491031478916e-05, + 3.495707896946e-05,  \
+ 3.500013339362e-05, + 3.503963205731e-05, + 3.507544985041e-05, + 3.510779701173e-05, + 3.513660522003e-05,  \
+ 3.516200173181e-05, + 3.518397639709e-05, + 3.520257494529e-05, + 3.521778013237e-05, + 3.522973274812e-05 ]

* Data table for Id-Vd at Vg = 0.54V
.param vd_data_vg0.54=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.54=[ \
+ 1.938900000000e-06, + 3.841400000000e-06, + 5.699500000000e-06, + 7.505700000000e-06, + 9.253200000000e-06,  \
+ 1.093630000000e-05, + 1.255020000000e-05, + 1.409140000000e-05, + 1.555710000000e-05, + 1.694560000000e-05,  \
+ 1.825610000000e-05, + 1.948900000000e-05, + 2.064520000000e-05, + 2.172660000000e-05, + 2.273560000000e-05,  \
+ 2.367520000000e-05, + 2.454860000000e-05, + 2.535910000000e-05, + 2.611000000000e-05, + 2.680480000000e-05,  \
+ 2.744660000000e-05, + 2.803870000000e-05, + 2.858420000000e-05, + 2.908620000000e-05, + 2.954800000000e-05,  \
+ 2.997260000000e-05, + 3.036320000000e-05, + 3.072260000000e-05, + 3.105380000000e-05, + 3.135940000000e-05,  \
+ 3.164190000000e-05, + 3.190350000000e-05, + 3.214640000000e-05, + 3.237250000000e-05, + 3.258350000000e-05,  \
+ 3.278100000000e-05, + 3.296620000000e-05, + 3.314050000000e-05, + 3.330490000000e-05, + 3.346040000000e-05,  \
+ 3.360790000000e-05, + 3.374810000000e-05, + 3.388170000000e-05, + 3.400930000000e-05, + 3.413150000000e-05,  \
+ 3.424870000000e-05, + 3.436140000000e-05, + 3.446990000000e-05, + 3.457460000000e-05, + 3.467580000000e-05,  \
+ 3.477370000000e-05, + 3.486870000000e-05, + 3.496100000000e-05, + 3.505060000000e-05, + 3.513800000000e-05,  \
+ 3.522310000000e-05, + 3.530620000000e-05, + 3.538730000000e-05, + 3.546670000000e-05, + 3.554440000000e-05,  \
+ 3.562050000000e-05, + 3.569520000000e-05, + 3.576850000000e-05, + 3.584040000000e-05, + 3.591120000000e-05,  \
+ 3.598080000000e-05, + 3.604930000000e-05, + 3.611670000000e-05, + 3.618320000000e-05, + 3.624870000000e-05,  \
+ 3.631340000000e-05, + 3.637720000000e-05, + 3.644020000000e-05, + 3.650250000000e-05, + 3.656400000000e-05,  \
+ 3.662480000000e-05, + 3.668500000000e-05, + 3.674450000000e-05, + 3.680340000000e-05, + 3.686170000000e-05 ]

.param id_pred_data_vg0.54=[ \
+ 1.982726535061e-06, + 3.902113239747e-06, + 5.756525642937e-06, + 7.544505642727e-06, + 9.264804975828e-06,  \
+ 1.091634796467e-05, + 1.249832013855e-05, + 1.401007291861e-05, + 1.545129198348e-05, + 1.682185393292e-05,  \
+ 1.812189366319e-05, + 1.935186737683e-05, + 2.051242146990e-05, + 2.160452364478e-05, + 2.262947964482e-05,  \
+ 2.358866855502e-05, + 2.448387240293e-05, + 2.531704871217e-05, + 2.609036440845e-05, + 2.680627512746e-05,  \
+ 2.746729238424e-05, + 2.807615790516e-05, + 2.863570000045e-05, + 2.914887503721e-05, + 2.961871905427e-05,  \
+ 3.004829675774e-05, + 3.044066514121e-05, + 3.079888178036e-05, + 3.112598722510e-05, + 3.142485729768e-05,  \
+ 3.169844960212e-05, + 3.194934688509e-05, + 3.218020079657e-05, + 3.239346464397e-05, + 3.259136756242e-05,  \
+ 3.277605457697e-05, + 3.294927046227e-05, + 3.311284497613e-05, + 3.326823512907e-05, + 3.341675328556e-05,  \
+ 3.355954606377e-05, + 3.369751604623e-05, + 3.383154944459e-05, + 3.396218875423e-05, + 3.408995980863e-05,  \
+ 3.421524394071e-05, + 3.433828227571e-05, + 3.445913898759e-05, + 3.457797392912e-05, + 3.469467992545e-05,  \
+ 3.480926789052e-05, + 3.492159914458e-05, + 3.503152373014e-05, + 3.513876770739e-05, + 3.524332314555e-05,  \
+ 3.534489893354e-05, + 3.544337501808e-05, + 3.553853413905e-05, + 3.563022492017e-05, + 3.571829074644e-05,  \
+ 3.580263681215e-05, + 3.588311607018e-05, + 3.595970112656e-05, + 3.603231860325e-05, + 3.610087951529e-05,  \
+ 3.616535570472e-05, + 3.622581185482e-05, + 3.628215767094e-05, + 3.633451244241e-05, + 3.638280250016e-05,  \
+ 3.642712596047e-05, + 3.646750235930e-05, + 3.650401718915e-05, + 3.653673906229e-05, + 3.656563785626e-05,  \
+ 3.659088062705e-05, + 3.661242019007e-05, + 3.663037910883e-05, + 3.664480322186e-05, + 3.665566619020e-05 ]

* Data table for Id-Vd at Vg = 0.55V
.param vd_data_vg0.55=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.55=[ \
+ 1.966800000000e-06, + 3.898700000000e-06, + 5.787600000000e-06, + 7.626000000000e-06, + 9.407200000000e-06,  \
+ 1.112540000000e-05, + 1.277610000000e-05, + 1.435530000000e-05, + 1.586030000000e-05, + 1.728930000000e-05,  \
+ 1.864140000000e-05, + 1.991650000000e-05, + 2.111550000000e-05, + 2.223980000000e-05, + 2.329160000000e-05,  \
+ 2.427360000000e-05, + 2.518890000000e-05, + 2.604060000000e-05, + 2.683190000000e-05, + 2.756610000000e-05,  \
+ 2.824640000000e-05, + 2.887580000000e-05, + 2.945740000000e-05, + 2.999430000000e-05, + 3.048940000000e-05,  \
+ 3.094590000000e-05, + 3.136660000000e-05, + 3.175450000000e-05, + 3.211240000000e-05, + 3.244300000000e-05,  \
+ 3.274880000000e-05, + 3.303220000000e-05, + 3.329530000000e-05, + 3.354010000000e-05, + 3.376850000000e-05,  \
+ 3.398210000000e-05, + 3.418220000000e-05, + 3.437040000000e-05, + 3.454760000000e-05, + 3.471510000000e-05,  \
+ 3.487370000000e-05, + 3.502420000000e-05, + 3.516750000000e-05, + 3.530410000000e-05, + 3.543480000000e-05,  \
+ 3.555990000000e-05, + 3.568000000000e-05, + 3.579550000000e-05, + 3.590670000000e-05, + 3.601410000000e-05,  \
+ 3.611800000000e-05, + 3.621850000000e-05, + 3.631600000000e-05, + 3.641070000000e-05, + 3.650280000000e-05,  \
+ 3.659240000000e-05, + 3.667980000000e-05, + 3.676510000000e-05, + 3.684840000000e-05, + 3.692980000000e-05,  \
+ 3.700960000000e-05, + 3.708770000000e-05, + 3.716430000000e-05, + 3.723950000000e-05, + 3.731330000000e-05,  \
+ 3.738590000000e-05, + 3.745720000000e-05, + 3.752740000000e-05, + 3.759660000000e-05, + 3.766470000000e-05,  \
+ 3.773190000000e-05, + 3.779810000000e-05, + 3.786350000000e-05, + 3.792800000000e-05, + 3.799180000000e-05,  \
+ 3.805470000000e-05, + 3.811700000000e-05, + 3.817860000000e-05, + 3.823950000000e-05, + 3.829980000000e-05 ]

.param id_pred_data_vg0.55=[ \
+ 2.010194730246e-06, + 3.959187888540e-06, + 5.845231935382e-06, + 7.666771416552e-06, + 9.422370203538e-06,  \
+ 1.111084478907e-05, + 1.273117377423e-05, + 1.428260933608e-05, + 1.576459442731e-05, + 1.717678242130e-05,  \
+ 1.851922206697e-05, + 1.979206921533e-05, + 2.099577468471e-05, + 2.213116560597e-05, + 2.319924169569e-05,  \
+ 2.420124597847e-05, + 2.513872372219e-05, + 2.601343032438e-05, + 2.682742735487e-05, + 2.758284099400e-05,  \
+ 2.828220371157e-05, + 2.892796648666e-05, + 2.952297727461e-05, + 3.007000079378e-05, + 3.057206413359e-05,  \
+ 3.103209703113e-05, + 3.145314534777e-05, + 3.183830209309e-05, + 3.219056583475e-05, + 3.251289599575e-05,  \
+ 3.280822376837e-05, + 3.307929029688e-05, + 3.332876753120e-05, + 3.355917579029e-05, + 3.377289649507e-05,  \
+ 3.397208667593e-05, + 3.415875486098e-05, + 3.433475169004e-05, + 3.450163654634e-05, + 3.466091293376e-05,  \
+ 3.481370396912e-05, + 3.496113160509e-05, + 3.510414200719e-05, + 3.524322470184e-05, + 3.537915545166e-05,  \
+ 3.551229383447e-05, + 3.564291837392e-05, + 3.577123163268e-05, + 3.589726191422e-05, + 3.602109791245e-05,  \
+ 3.614255103457e-05, + 3.626171033829e-05, + 3.637824454927e-05, + 3.649201156804e-05, + 3.660289876279e-05,  \
+ 3.671063459478e-05, + 3.681501846586e-05, + 3.691587160574e-05, + 3.701302004629e-05, + 3.710630990099e-05,  \
+ 3.719556360011e-05, + 3.728063260496e-05, + 3.736155347724e-05, + 3.743810812011e-05, + 3.751027506951e-05,  \
+ 3.757805650821e-05, + 3.764148281334e-05, + 3.770039198571e-05, + 3.775489960390e-05, + 3.780511360674e-05,  \
+ 3.785099055676e-05, + 3.789258567849e-05, + 3.792994473770e-05, + 3.796322322160e-05, + 3.799241676461e-05,  \
+ 3.801766652032e-05, + 3.803895633610e-05, + 3.805641827057e-05, + 3.807006167335e-05, + 3.808014735114e-05 ]

* Data table for Id-Vd at Vg = 0.56V
.param vd_data_vg0.56=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.56=[ \
+ 1.993600000000e-06, + 3.953400000000e-06, + 5.871700000000e-06, + 7.740800000000e-06, + 9.554300000000e-06,  \
+ 1.130630000000e-05, + 1.299200000000e-05, + 1.460770000000e-05, + 1.615050000000e-05, + 1.761850000000e-05,  \
+ 1.901060000000e-05, + 2.032660000000e-05, + 2.156690000000e-05, + 2.273290000000e-05, + 2.382650000000e-05,  \
+ 2.485000000000e-05, + 2.580630000000e-05, + 2.669850000000e-05, + 2.752950000000e-05, + 2.830270000000e-05,  \
+ 2.902090000000e-05, + 2.968740000000e-05, + 3.030500000000e-05, + 3.087670000000e-05, + 3.140530000000e-05,  \
+ 3.189390000000e-05, + 3.234520000000e-05, + 3.276220000000e-05, + 3.314760000000e-05, + 3.350400000000e-05,  \
+ 3.383400000000e-05, + 3.413990000000e-05, + 3.442410000000e-05, + 3.468860000000e-05, + 3.493520000000e-05,  \
+ 3.516570000000e-05, + 3.538160000000e-05, + 3.558440000000e-05, + 3.577530000000e-05, + 3.595540000000e-05,  \
+ 3.612570000000e-05, + 3.628730000000e-05, + 3.644080000000e-05, + 3.658700000000e-05, + 3.672660000000e-05,  \
+ 3.686010000000e-05, + 3.698800000000e-05, + 3.711090000000e-05, + 3.722920000000e-05, + 3.734320000000e-05,  \
+ 3.745320000000e-05, + 3.755960000000e-05, + 3.766270000000e-05, + 3.776260000000e-05, + 3.785970000000e-05,  \
+ 3.795410000000e-05, + 3.804600000000e-05, + 3.813560000000e-05, + 3.822300000000e-05, + 3.830840000000e-05,  \
+ 3.839200000000e-05, + 3.847370000000e-05, + 3.855380000000e-05, + 3.863230000000e-05, + 3.870930000000e-05,  \
+ 3.878500000000e-05, + 3.885930000000e-05, + 3.893240000000e-05, + 3.900430000000e-05, + 3.907510000000e-05,  \
+ 3.914490000000e-05, + 3.921360000000e-05, + 3.928140000000e-05, + 3.934830000000e-05, + 3.941440000000e-05,  \
+ 3.947960000000e-05, + 3.954400000000e-05, + 3.960770000000e-05, + 3.967060000000e-05, + 3.973290000000e-05 ]

.param id_pred_data_vg0.56=[ \
+ 2.036487130681e-06, + 4.013780853711e-06, + 5.930037586950e-06, + 7.783600012772e-06, + 9.572932322044e-06,  \
+ 1.129670214141e-05, + 1.295377893257e-05, + 1.454325392842e-05, + 1.606436664588e-05, + 1.751671661623e-05,  \
+ 1.890002953587e-05, + 2.021435124334e-05, + 2.145996259060e-05, + 2.263745933305e-05, + 2.374762771069e-05,  \
+ 2.479154150933e-05, + 2.577055856818e-05, + 2.668622735655e-05, + 2.754039174761e-05, + 2.833511098288e-05,  \
+ 2.907264643000e-05, + 2.975532261189e-05, + 3.038592229132e-05, + 3.096709144302e-05, + 3.150167322019e-05,  \
+ 3.199262311682e-05, + 3.244288047426e-05, + 3.285559971118e-05, + 3.323369601276e-05, + 3.358014364494e-05,  \
+ 3.389793033421e-05, + 3.418983658776e-05, + 3.445859634667e-05, + 3.470687501249e-05, + 3.493703225104e-05,  \
+ 3.515143616823e-05, + 3.535213778378e-05, + 3.554102586349e-05, + 3.571987086616e-05, + 3.589031693991e-05,  \
+ 3.605350997532e-05, + 3.621078169090e-05, + 3.636299661594e-05, + 3.651092993096e-05, + 3.665524782264e-05,  \
+ 3.679655506858e-05, + 3.693500417285e-05, + 3.707094001584e-05, + 3.720442102349e-05, + 3.733551056939e-05,  \
+ 3.746421585674e-05, + 3.759034996619e-05, + 3.771378222154e-05, + 3.783435633522e-05, + 3.795185766649e-05,  \
+ 3.806606575381e-05, + 3.817667522526e-05, + 3.828359156614e-05, + 3.838657059532e-05, + 3.848537744489e-05,  \
+ 3.857997544401e-05, + 3.867005172651e-05, + 3.875565453200e-05, + 3.883654484525e-05, + 3.891274445778e-05,  \
+ 3.898417598975e-05, + 3.905087003659e-05, + 3.911273117410e-05, + 3.916983961972e-05, + 3.922227297153e-05,  \
+ 3.927001984266e-05, + 3.931313491194e-05, + 3.935163374990e-05, + 3.938581998227e-05, + 3.941554496123e-05,  \
+ 3.944091062294e-05, + 3.946217300836e-05, + 3.947934455937e-05, + 3.949248060962e-05, + 3.950170066673e-05 ]

* Data table for Id-Vd at Vg = 0.57V
.param vd_data_vg0.57=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.57=[ \
+ 2.019100000000e-06, + 4.005700000000e-06, + 5.952000000000e-06, + 7.850600000000e-06, + 9.694900000000e-06,  \
+ 1.147910000000e-05, + 1.319850000000e-05, + 1.484920000000e-05, + 1.642830000000e-05, + 1.793380000000e-05,  \
+ 1.936450000000e-05, + 2.071980000000e-05, + 2.200020000000e-05, + 2.320660000000e-05, + 2.434070000000e-05,  \
+ 2.540480000000e-05, + 2.640120000000e-05, + 2.733300000000e-05, + 2.820320000000e-05, + 2.901460000000e-05,  \
+ 2.977040000000e-05, + 3.047350000000e-05, + 3.112680000000e-05, + 3.173320000000e-05, + 3.229530000000e-05,  \
+ 3.281620000000e-05, + 3.329840000000e-05, + 3.374490000000e-05, + 3.415820000000e-05, + 3.454110000000e-05,  \
+ 3.489600000000e-05, + 3.522540000000e-05, + 3.553150000000e-05, + 3.581640000000e-05, + 3.608200000000e-05,  \
+ 3.633030000000e-05, + 3.656280000000e-05, + 3.678090000000e-05, + 3.698610000000e-05, + 3.717960000000e-05,  \
+ 3.736240000000e-05, + 3.753550000000e-05, + 3.769990000000e-05, + 3.785620000000e-05, + 3.800520000000e-05,  \
+ 3.814760000000e-05, + 3.828390000000e-05, + 3.841470000000e-05, + 3.854030000000e-05, + 3.866120000000e-05,  \
+ 3.877780000000e-05, + 3.889040000000e-05, + 3.899930000000e-05, + 3.910480000000e-05, + 3.920710000000e-05,  \
+ 3.930650000000e-05, + 3.940320000000e-05, + 3.949730000000e-05, + 3.958910000000e-05, + 3.967860000000e-05,  \
+ 3.976610000000e-05, + 3.985170000000e-05, + 3.993540000000e-05, + 4.001740000000e-05, + 4.009780000000e-05,  \
+ 4.017660000000e-05, + 4.025410000000e-05, + 4.033010000000e-05, + 4.040490000000e-05, + 4.047850000000e-05,  \
+ 4.055100000000e-05, + 4.062230000000e-05, + 4.069260000000e-05, + 4.076200000000e-05, + 4.083030000000e-05,  \
+ 4.089780000000e-05, + 4.096450000000e-05, + 4.103030000000e-05, + 4.109540000000e-05, + 4.115970000000e-05 ]

.param id_pred_data_vg0.57=[ \
+ 2.061634586425e-06, + 4.065953544341e-06, + 6.011049990775e-06, + 7.895150920376e-06, + 9.716676140670e-06,  \
+ 1.147417235188e-05, + 1.316638212302e-05, + 1.479228143580e-05, + 1.635095963138e-05, + 1.784185878932e-05,  \
+ 1.926462180563e-05, + 2.061900158878e-05, + 2.190518760472e-05, + 2.312358206837e-05, + 2.427480794722e-05,  \
+ 2.535963896662e-05, + 2.637937446707e-05, + 2.733530884143e-05, + 2.822916911100e-05, + 2.906274457928e-05,  \
+ 2.983824771945e-05, + 3.055778128328e-05, + 3.122402296867e-05, + 3.183943452314e-05, + 3.240680962335e-05,  \
+ 3.292906912975e-05, + 3.340904149809e-05, + 3.384983341675e-05, + 3.425429742492e-05, + 3.462551321718e-05,  \
+ 3.496639641526e-05, + 3.527981461957e-05, + 3.556850351742e-05, + 3.583523634006e-05, + 3.608251172409e-05,  \
+ 3.631267027231e-05, + 3.652787396277e-05, + 3.673025741591e-05, + 3.692163561936e-05, + 3.710358578246e-05,  \
+ 3.727762763447e-05, + 3.744502391783e-05, + 3.760676481761e-05, + 3.776375815505e-05, + 3.791678645939e-05,  \
+ 3.806640437688e-05, + 3.821291189524e-05, + 3.835669602267e-05, + 3.849781838653e-05, + 3.863644815283e-05,  \
+ 3.877252573147e-05, + 3.890591760864e-05, + 3.903646313120e-05, + 3.916406931239e-05, + 3.928847108909e-05,  \
+ 3.940933442209e-05, + 3.952659513743e-05, + 3.963990049670e-05, + 3.974907143856e-05, + 3.985385410488e-05,  \
+ 3.995406150352e-05, + 4.004952614196e-05, + 4.014024409116e-05, + 4.022583365440e-05, + 4.030648342450e-05,  \
+ 4.038201659569e-05, + 4.045233556099e-05, + 4.051761425217e-05, + 4.057770587679e-05, + 4.063268133905e-05,  \
+ 4.068260979693e-05, + 4.072758631082e-05, + 4.076766606886e-05, + 4.080296523171e-05, + 4.083344811079e-05,  \
+ 4.085937704076e-05, + 4.088081524969e-05, + 4.089790374564e-05, + 4.091061440704e-05, + 4.091919108760e-05 ]

* Data table for Id-Vd at Vg = 0.58V
.param vd_data_vg0.58=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.58=[ \
+ 2.043500000000e-06, + 4.055600000000e-06, + 6.028800000000e-06, + 7.955500000000e-06, + 9.829200000000e-06,  \
+ 1.164430000000e-05, + 1.339590000000e-05, + 1.508020000000e-05, + 1.669420000000e-05, + 1.823570000000e-05,  \
+ 1.970340000000e-05, + 2.109680000000e-05, + 2.241580000000e-05, + 2.366140000000e-05, + 2.483500000000e-05,  \
+ 2.593850000000e-05, + 2.697420000000e-05, + 2.794480000000e-05, + 2.885320000000e-05, + 2.970230000000e-05,  \
+ 3.049510000000e-05, + 3.123430000000e-05, + 3.192300000000e-05, + 3.256370000000e-05, + 3.315930000000e-05,  \
+ 3.371240000000e-05, + 3.422570000000e-05, + 3.470190000000e-05, + 3.514360000000e-05, + 3.555350000000e-05,  \
+ 3.593390000000e-05, + 3.628730000000e-05, + 3.661600000000e-05, + 3.692210000000e-05, + 3.720760000000e-05,  \
+ 3.747440000000e-05, + 3.772410000000e-05, + 3.795840000000e-05, + 3.817870000000e-05, + 3.838620000000e-05,  \
+ 3.858210000000e-05, + 3.876740000000e-05, + 3.894320000000e-05, + 3.911020000000e-05, + 3.926930000000e-05,  \
+ 3.942100000000e-05, + 3.956610000000e-05, + 3.970510000000e-05, + 3.983850000000e-05, + 3.996670000000e-05,  \
+ 4.009020000000e-05, + 4.020930000000e-05, + 4.032440000000e-05, + 4.043570000000e-05, + 4.054360000000e-05,  \
+ 4.064820000000e-05, + 4.074990000000e-05, + 4.084880000000e-05, + 4.094510000000e-05, + 4.103900000000e-05,  \
+ 4.113060000000e-05, + 4.122010000000e-05, + 4.130760000000e-05, + 4.139330000000e-05, + 4.147710000000e-05,  \
+ 4.155930000000e-05, + 4.164000000000e-05, + 4.171920000000e-05, + 4.179700000000e-05, + 4.187350000000e-05,  \
+ 4.194870000000e-05, + 4.202270000000e-05, + 4.209560000000e-05, + 4.216750000000e-05, + 4.223830000000e-05,  \
+ 4.230820000000e-05, + 4.237710000000e-05, + 4.244520000000e-05, + 4.251240000000e-05, + 4.257880000000e-05 ]

.param id_pred_data_vg0.58=[ \
+ 2.085659943987e-06, + 4.115761548746e-06, + 6.088336376706e-06, + 8.001574897207e-06, + 9.853797382675e-06,  \
+ 1.164347719168e-05, + 1.336925939540e-05, + 1.503001200035e-05, + 1.662467591814e-05, + 1.815264695324e-05,  \
+ 1.961328380276e-05, + 2.100637299009e-05, + 2.233179780887e-05, + 2.358984347666e-05, + 2.478086753399e-05,  \
+ 2.590570133179e-05, + 2.696526047657e-05, + 2.796073764330e-05, + 2.889364332077e-05, + 2.976565447170e-05,  \
+ 3.057868976612e-05, + 3.133499034448e-05, + 3.203671367373e-05, + 3.268646774814e-05, + 3.328686943860e-05,  \
+ 3.384067269508e-05, + 3.435079546762e-05, + 3.482004976831e-05, + 3.525139945850e-05, + 3.564793296391e-05,  \
+ 3.601251453802e-05, + 3.634799504653e-05, + 3.665727410407e-05, + 3.694316386827e-05, + 3.720805143530e-05,  \
+ 3.745453432202e-05, + 3.768491078517e-05, + 3.790122704231e-05, + 3.810546375462e-05, + 3.829941852018e-05,  \
+ 3.848472049867e-05, + 3.866255341563e-05, + 3.883414508891e-05, + 3.900053765392e-05, + 3.916242567357e-05,  \
+ 3.932059669751e-05, + 3.947535573388e-05, + 3.962710266933e-05, + 3.977612417657e-05, + 3.992244091933e-05,  \
+ 4.006602604932e-05, + 4.020685824798e-05, + 4.034481033159e-05, + 4.047962604091e-05, + 4.061119034304e-05,  \
+ 4.073911230080e-05, + 4.086313587322e-05, + 4.098312725546e-05, + 4.109877969313e-05, + 4.120987141505e-05,  \
+ 4.131608860916e-05, + 4.141741155763e-05, + 4.151357112278e-05, + 4.160438198596e-05, + 4.168982959527e-05,  \
+ 4.176986636594e-05, + 4.184431454632e-05, + 4.191327985609e-05, + 4.197676131298e-05, + 4.203471653454e-05,  \
+ 4.208729071252e-05, + 4.213446256472e-05, + 4.217636858812e-05, + 4.221308947308e-05, + 4.224486838211e-05,  \
+ 4.227156998240e-05, + 4.229342921462e-05, + 4.231062310282e-05, + 4.232320712617e-05, + 4.233135550749e-05 ]

* Data table for Id-Vd at Vg = 0.59V
.param vd_data_vg0.59=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.59=[ \
+ 2.066800000000e-06, + 4.103400000000e-06, + 6.102100000000e-06, + 8.055700000000e-06, + 9.957700000000e-06,  \
+ 1.180230000000e-05, + 1.358480000000e-05, + 1.530130000000e-05, + 1.694870000000e-05, + 1.852480000000e-05,  \
+ 2.002820000000e-05, + 2.145810000000e-05, + 2.281460000000e-05, + 2.409810000000e-05, + 2.530990000000e-05,  \
+ 2.645170000000e-05, + 2.752560000000e-05, + 2.853420000000e-05, + 2.948010000000e-05, + 3.036620000000e-05,  \
+ 3.119520000000e-05, + 3.197010000000e-05, + 3.269360000000e-05, + 3.336830000000e-05, + 3.399700000000e-05,  \
+ 3.458230000000e-05, + 3.512670000000e-05, + 3.563280000000e-05, + 3.610320000000e-05, + 3.654030000000e-05,  \
+ 3.694670000000e-05, + 3.732470000000e-05, + 3.767660000000e-05, + 3.800460000000e-05, + 3.831060000000e-05,  \
+ 3.859660000000e-05, + 3.886440000000e-05, + 3.911550000000e-05, + 3.935150000000e-05, + 3.957370000000e-05,  \
+ 3.978330000000e-05, + 3.998150000000e-05, + 4.016920000000e-05, + 4.034750000000e-05, + 4.051710000000e-05,  \
+ 4.067870000000e-05, + 4.083300000000e-05, + 4.098070000000e-05, + 4.112220000000e-05, + 4.125820000000e-05,  \
+ 4.138890000000e-05, + 4.151490000000e-05, + 4.163640000000e-05, + 4.175390000000e-05, + 4.186760000000e-05,  \
+ 4.197780000000e-05, + 4.208470000000e-05, + 4.218860000000e-05, + 4.228970000000e-05, + 4.238810000000e-05,  \
+ 4.248400000000e-05, + 4.257770000000e-05, + 4.266910000000e-05, + 4.275850000000e-05, + 4.284610000000e-05,  \
+ 4.293180000000e-05, + 4.301580000000e-05, + 4.309820000000e-05, + 4.317910000000e-05, + 4.325860000000e-05,  \
+ 4.333670000000e-05, + 4.341350000000e-05, + 4.348910000000e-05, + 4.356360000000e-05, + 4.363690000000e-05,  \
+ 4.370920000000e-05, + 4.378050000000e-05, + 4.385090000000e-05, + 4.392030000000e-05, + 4.398890000000e-05 ]

.param id_pred_data_vg0.59=[ \
+ 2.108589542331e-06, + 4.163260164205e-06, + 6.162013305584e-06, + 8.103001164272e-06, + 9.984461212298e-06,  \
+ 1.180481660413e-05, + 1.356264605420e-05, + 1.525667263195e-05, + 1.688583244686e-05, + 1.844930957304e-05,  \
+ 1.994642530917e-05, + 2.137670817319e-05, + 2.274006939842e-05, + 2.403644524748e-05, + 2.526622774894e-05,  \
+ 2.642992418259e-05, + 2.752837739536e-05, + 2.856256352970e-05, + 2.953385032015e-05, + 3.044375916943e-05,  \
+ 3.129399396130e-05, + 3.208658163203e-05, + 3.282376012066e-05, + 3.350781393237e-05, + 3.414130333113e-05,  \
+ 3.472686628811e-05, + 3.526726621203e-05, + 3.576543997042e-05, + 3.622417920269e-05, + 3.664651012514e-05,  \
+ 3.703528775077e-05, + 3.739348612726e-05, + 3.772396448767e-05, + 3.802941326285e-05, + 3.831257672573e-05,  \
+ 3.857597534079e-05, + 3.882195065671e-05, + 3.905272373231e-05, + 3.927035642846e-05, + 3.947679069825e-05,  \
+ 3.967357741203e-05, + 3.986218755017e-05, + 4.004391412309e-05, + 4.021986300359e-05, + 4.039093437314e-05,  \
+ 4.055777986650e-05, + 4.072101910424e-05, + 4.088094807230e-05, + 4.103797291464e-05, + 4.119207005715e-05,  \
+ 4.134337723372e-05, + 4.149182874244e-05, + 4.163728131971e-05, + 4.177956492640e-05, + 4.191839470877e-05,  \
+ 4.205356177408e-05, + 4.218476293318e-05, + 4.231174418237e-05, + 4.243421863066e-05, + 4.255188396201e-05,  \
+ 4.266452997399e-05, + 4.277193511371e-05, + 4.287393501727e-05, + 4.297039005905e-05, + 4.306110640755e-05,  \
+ 4.314595091273e-05, + 4.322504471929e-05, + 4.329818184488e-05, + 4.336545462138e-05, + 4.342682004790e-05,  \
+ 4.348233458586e-05, + 4.353219468612e-05, + 4.357640282251e-05, + 4.361496779893e-05, + 4.364813321445e-05,  \
+ 4.367601577542e-05, + 4.369868431240e-05, + 4.371628245281e-05, + 4.372903444164e-05, + 4.373699193820e-05 ]

* Data table for Id-Vd at Vg = 0.60V
.param vd_data_vg0.60=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.60=[ \
+ 2.089000000000e-06, + 4.149000000000e-06, + 6.172200000000e-06, + 8.151600000000e-06, + 1.008050000000e-05,  \
+ 1.195340000000e-05, + 1.376550000000e-05, + 1.551280000000e-05, + 1.719230000000e-05, + 1.880170000000e-05,  \
+ 2.033940000000e-05, + 2.180460000000e-05, + 2.319700000000e-05, + 2.451710000000e-05, + 2.576600000000e-05,  \
+ 2.694500000000e-05, + 2.805610000000e-05, + 2.910170000000e-05, + 3.008430000000e-05, + 3.100660000000e-05,  \
+ 3.187130000000e-05, + 3.268110000000e-05, + 3.343890000000e-05, + 3.414720000000e-05, + 3.480870000000e-05,  \
+ 3.542580000000e-05, + 3.600120000000e-05, + 3.653720000000e-05, + 3.703630000000e-05, + 3.750110000000e-05,  \
+ 3.793380000000e-05, + 3.833680000000e-05, + 3.871240000000e-05, + 3.906280000000e-05, + 3.938990000000e-05,  \
+ 3.969580000000e-05, + 3.998220000000e-05, + 4.025080000000e-05, + 4.050320000000e-05, + 4.074070000000e-05,  \
+ 4.096460000000e-05, + 4.117630000000e-05, + 4.137660000000e-05, + 4.156660000000e-05, + 4.174720000000e-05,  \
+ 4.191920000000e-05, + 4.208320000000e-05, + 4.224000000000e-05, + 4.239020000000e-05, + 4.253420000000e-05,  \
+ 4.267260000000e-05, + 4.280570000000e-05, + 4.293410000000e-05, + 4.305800000000e-05, + 4.317780000000e-05,  \
+ 4.329380000000e-05, + 4.340620000000e-05, + 4.351530000000e-05, + 4.362130000000e-05, + 4.372450000000e-05,  \
+ 4.382490000000e-05, + 4.392290000000e-05, + 4.401850000000e-05, + 4.411190000000e-05, + 4.420320000000e-05,  \
+ 4.429250000000e-05, + 4.438000000000e-05, + 4.446580000000e-05, + 4.454990000000e-05, + 4.463250000000e-05,  \
+ 4.471360000000e-05, + 4.479330000000e-05, + 4.487170000000e-05, + 4.494880000000e-05, + 4.502480000000e-05,  \
+ 4.509960000000e-05, + 4.517330000000e-05, + 4.524610000000e-05, + 4.531780000000e-05, + 4.538860000000e-05 ]

.param id_pred_data_vg0.60=[ \
+ 2.130443899659e-06, + 4.208500904497e-06, + 6.232170271687e-06, + 8.199548465200e-06, + 1.010882406263e-05,  \
+ 1.195842021843e-05, + 1.374678962748e-05, + 1.547260791995e-05, + 1.713474353892e-05, + 1.873221481219e-05,  \
+ 2.026430243859e-05, + 2.173043321818e-05, + 2.313031262020e-05, + 2.446379279718e-05, + 2.573106758064e-05,  \
+ 2.693257993087e-05, + 2.806883654557e-05, + 2.914091222920e-05, + 3.014980393345e-05, + 3.109695098829e-05,  \
+ 3.198390666512e-05, + 3.281255194452e-05, + 3.358485104400e-05, + 3.430308192037e-05, + 3.496967838146e-05,  \
+ 3.558716183761e-05, + 3.615811583586e-05, + 3.668538469356e-05, + 3.717183906701e-05, + 3.762042179005e-05,  \
+ 3.803389729001e-05, + 3.841530531645e-05, + 3.876741735439e-05, + 3.909309642040e-05, + 3.939510970667e-05,  \
+ 3.967590106186e-05, + 3.993799211457e-05, + 4.018371619168e-05, + 4.041528074595e-05, + 4.063439846504e-05,  \
+ 4.084311251063e-05, + 4.104287509108e-05, + 4.123502068978e-05, + 4.142082500039e-05, + 4.160116659477e-05,  \
+ 4.177695984254e-05, + 4.194874614768e-05, + 4.211702733301e-05, + 4.228206686093e-05, + 4.244423689670e-05,  \
+ 4.260339555913e-05, + 4.275958810467e-05, + 4.291263823688e-05, + 4.306256581913e-05, + 4.320883163018e-05,  \
+ 4.335150937550e-05, + 4.349003720563e-05, + 4.362427425804e-05, + 4.375376127427e-05, + 4.387843364384e-05,  \
+ 4.399777892104e-05, + 4.411173897097e-05, + 4.421988269314e-05, + 4.432236775756e-05, + 4.441864912224e-05,  \
+ 4.450893044122e-05, + 4.459294417757e-05, + 4.467065533390e-05, + 4.474215165828e-05, + 4.480742572923e-05,  \
+ 4.486638019443e-05, + 4.491932108067e-05, + 4.496618596022e-05, + 4.500696610194e-05, + 4.504209118750e-05,  \
+ 4.507138175541e-05, + 4.509516031248e-05, + 4.511366445513e-05, + 4.512673982390e-05, + 4.513486637734e-05 ]

* Data table for Id-Vd at Vg = 0.61V
.param vd_data_vg0.61=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.61=[ \
+ 2.110400000000e-06, + 4.192600000000e-06, + 6.239300000000e-06, + 8.243200000000e-06, + 1.019800000000e-05,  \
+ 1.209800000000e-05, + 1.393840000000e-05, + 1.571530000000e-05, + 1.742560000000e-05, + 1.906680000000e-05,  \
+ 2.063750000000e-05, + 2.213660000000e-05, + 2.356380000000e-05, + 2.491930000000e-05, + 2.620390000000e-05,  \
+ 2.741900000000e-05, + 2.856630000000e-05, + 2.964800000000e-05, + 3.066640000000e-05, + 3.162400000000e-05,  \
+ 3.252360000000e-05, + 3.336780000000e-05, + 3.415930000000e-05, + 3.490070000000e-05, + 3.559450000000e-05,  \
+ 3.624320000000e-05, + 3.684920000000e-05, + 3.741490000000e-05, + 3.794280000000e-05, + 3.843520000000e-05,  \
+ 3.889450000000e-05, + 3.932290000000e-05, + 3.972260000000e-05, + 4.009580000000e-05, + 4.044460000000e-05,  \
+ 4.077090000000e-05, + 4.107650000000e-05, + 4.136320000000e-05, + 4.163250000000e-05, + 4.188590000000e-05,  \
+ 4.212480000000e-05, + 4.235040000000e-05, + 4.256390000000e-05, + 4.276620000000e-05, + 4.295830000000e-05,  \
+ 4.314110000000e-05, + 4.331530000000e-05, + 4.348170000000e-05, + 4.364090000000e-05, + 4.379330000000e-05,  \
+ 4.393970000000e-05, + 4.408040000000e-05, + 4.421590000000e-05, + 4.434660000000e-05, + 4.447280000000e-05,  \
+ 4.459480000000e-05, + 4.471290000000e-05, + 4.482750000000e-05, + 4.493870000000e-05, + 4.504690000000e-05,  \
+ 4.515200000000e-05, + 4.525450000000e-05, + 4.535440000000e-05, + 4.545190000000e-05, + 4.554710000000e-05,  \
+ 4.564030000000e-05, + 4.573140000000e-05, + 4.582060000000e-05, + 4.590810000000e-05, + 4.599390000000e-05,  \
+ 4.607810000000e-05, + 4.616080000000e-05, + 4.624210000000e-05, + 4.632200000000e-05, + 4.640060000000e-05,  \
+ 4.647810000000e-05, + 4.655430000000e-05, + 4.662950000000e-05, + 4.670360000000e-05, + 4.677660000000e-05 ]

.param id_pred_data_vg0.61=[ \
+ 2.151242224500e-06, + 4.251544014551e-06, + 6.298883672571e-06, + 8.291330304928e-06, + 1.022709620884e-05,  \
+ 1.210446003824e-05, + 1.392190402839e-05, + 1.567804836668e-05, + 1.737165934173e-05, + 1.900169008877e-05,  \
+ 2.056732977508e-05, + 2.206783974543e-05, + 2.350289825699e-05, + 2.487215708243e-05, + 2.617575810291e-05,  \
+ 2.741387579590e-05, + 2.858703621314e-05, + 2.969600376673e-05, + 3.074172811466e-05, + 3.172537835781e-05,  \
+ 3.264846760430e-05, + 3.351270279381e-05, + 3.431986930082e-05, + 3.507211105898e-05, + 3.577165625757e-05,  \
+ 3.642101451987e-05, + 3.702271176735e-05, + 3.757939091884e-05, + 3.809390007518e-05, + 3.856902185362e-05,  \
+ 3.900764844730e-05, + 3.941272851080e-05, + 3.978699642175e-05, + 4.013344645500e-05, + 4.045468522236e-05,  \
+ 4.075344448211e-05, + 4.103220060642e-05, + 4.129331689910e-05, + 4.153907895670e-05, + 4.177145892754e-05,  \
+ 4.199246068310e-05, + 4.220360147883e-05, + 4.240651993314e-05, + 4.260235436959e-05, + 4.279224813217e-05,  \
+ 4.297708903323e-05, + 4.315759644669e-05, + 4.333428572863e-05, + 4.350761810201e-05, + 4.367774090497e-05,  \
+ 4.384482308524e-05, + 4.400884616189e-05, + 4.416969335580e-05, + 4.432735178852e-05, + 4.448138861335e-05,  \
+ 4.463154939003e-05, + 4.477762740862e-05, + 4.491930798395e-05, + 4.505616270762e-05, + 4.518794885371e-05,  \
+ 4.531435748504e-05, + 4.543514951365e-05, + 4.555001607514e-05, + 4.565871320665e-05, + 4.576108622132e-05,  \
+ 4.585711460095e-05, + 4.594651632942e-05, + 4.602939909091e-05, + 4.610557472915e-05, + 4.617504382622e-05,  \
+ 4.623795524822e-05, + 4.629432514776e-05, + 4.634421486116e-05, + 4.638774640625e-05, + 4.642505882657e-05,  \
+ 4.645639884984e-05, + 4.648170870496e-05, + 4.650127084460e-05, + 4.651523402572e-05, + 4.652374482248e-05 ]

* Data table for Id-Vd at Vg = 0.62V
.param vd_data_vg0.62=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.62=[ \
+ 2.130700000000e-06, + 4.234400000000e-06, + 6.303500000000e-06, + 8.331000000000e-06, + 1.031050000000e-05,  \
+ 1.223640000000e-05, + 1.410390000000e-05, + 1.590920000000e-05, + 1.764890000000e-05, + 1.932080000000e-05,  \
+ 2.092320000000e-05, + 2.245490000000e-05, + 2.391550000000e-05, + 2.530510000000e-05, + 2.662440000000e-05,  \
+ 2.787440000000e-05, + 2.905690000000e-05, + 3.017360000000e-05, + 3.122680000000e-05, + 3.221900000000e-05,  \
+ 3.315280000000e-05, + 3.403060000000e-05, + 3.485520000000e-05, + 3.562900000000e-05, + 3.635460000000e-05,  \
+ 3.703440000000e-05, + 3.767080000000e-05, + 3.826610000000e-05, + 3.882260000000e-05, + 3.934260000000e-05,  \
+ 3.982850000000e-05, + 4.028240000000e-05, + 4.070650000000e-05, + 4.110290000000e-05, + 4.147380000000e-05,  \
+ 4.182090000000e-05, + 4.214630000000e-05, + 4.245150000000e-05, + 4.273830000000e-05, + 4.300820000000e-05,  \
+ 4.326260000000e-05, + 4.350270000000e-05, + 4.372980000000e-05, + 4.394490000000e-05, + 4.414910000000e-05,  \
+ 4.434320000000e-05, + 4.452800000000e-05, + 4.470440000000e-05, + 4.487300000000e-05, + 4.503430000000e-05,  \
+ 4.518900000000e-05, + 4.533760000000e-05, + 4.548060000000e-05, + 4.561830000000e-05, + 4.575120000000e-05,  \
+ 4.587950000000e-05, + 4.600370000000e-05, + 4.612400000000e-05, + 4.624060000000e-05, + 4.635390000000e-05,  \
+ 4.646400000000e-05, + 4.657110000000e-05, + 4.667550000000e-05, + 4.677730000000e-05, + 4.687660000000e-05,  \
+ 4.697370000000e-05, + 4.706860000000e-05, + 4.716150000000e-05, + 4.725240000000e-05, + 4.734150000000e-05,  \
+ 4.742900000000e-05, + 4.751470000000e-05, + 4.759900000000e-05, + 4.768180000000e-05, + 4.776320000000e-05,  \
+ 4.784330000000e-05, + 4.792220000000e-05, + 4.799980000000e-05, + 4.807630000000e-05, + 4.815180000000e-05 ]

.param id_pred_data_vg0.62=[ \
+ 2.171011292376e-06, + 4.292435187381e-06, + 6.362226413330e-06, + 8.378471829928e-06, + 1.033935404848e-05,  \
+ 1.224316132721e-05, + 1.408826836268e-05, + 1.587329781614e-05, + 1.759692691849e-05, + 1.925804681377e-05,  \
+ 2.085580345010e-05, + 2.238929271698e-05, + 2.385817628237e-05, + 2.526193333324e-05, + 2.660059835762e-05,  \
+ 2.787424949929e-05, + 2.908316688263e-05, + 3.022809483809e-05, + 3.130975004751e-05, + 3.232926828787e-05,  \
+ 3.328779595904e-05, + 3.418714302825e-05, + 3.502872452373e-05, + 3.581470227800e-05, + 3.654717875179e-05,  \
+ 3.722832596395e-05, + 3.786075933021e-05, + 3.844690450933e-05, + 3.898972077877e-05, + 3.949175588787e-05,  \
+ 3.995584876975e-05, + 4.038502462208e-05, + 4.078198136995e-05, + 4.114960989682e-05, + 4.149061314820e-05,  \
+ 4.180778574664e-05, + 4.210367158521e-05, + 4.238065768732e-05, + 4.264106719347e-05, + 4.288709606044e-05,  \
+ 4.312066135753e-05, + 4.334363329690e-05, + 4.355747325462e-05, + 4.376363154734e-05, + 4.396322947287e-05,  \
+ 4.415734074428e-05, + 4.434669455804e-05, + 4.453194444068e-05, + 4.471356776776e-05, + 4.489178536460e-05,  \
+ 4.506682118517e-05, + 4.523882351350e-05, + 4.540745947452e-05, + 4.557283842587e-05, + 4.573464902933e-05,  \
+ 4.589254094753e-05, + 4.604638888850e-05, + 4.619569750503e-05, + 4.634010932932e-05, + 4.647937312257e-05,  \
+ 4.661304068577e-05, + 4.674099385738e-05, + 4.686278123700e-05, + 4.697815515101e-05, + 4.708711712738e-05,  \
+ 4.718921161839e-05, + 4.728450832772e-05, + 4.737273586215e-05, + 4.745408215967e-05, + 4.752829918289e-05,  \
+ 4.759555129567e-05, + 4.765585006680e-05, + 4.770939005539e-05, + 4.775602996233e-05, + 4.779599112226e-05,  \
+ 4.782962379977e-05, + 4.785682242073e-05, + 4.787792116986e-05, + 4.789302831341e-05, + 4.790238454007e-05 ]

* Data table for Id-Vd at Vg = 0.63V
.param vd_data_vg0.63=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.63=[ \
+ 2.150300000000e-06, + 4.274300000000e-06, + 6.364900000000e-06, + 8.414900000000e-06, + 1.041810000000e-05,  \
+ 1.236890000000e-05, + 1.426240000000e-05, + 1.609480000000e-05, + 1.786290000000e-05, + 1.956420000000e-05,  \
+ 2.119690000000e-05, + 2.276000000000e-05, + 2.425280000000e-05, + 2.567520000000e-05, + 2.702790000000e-05,  \
+ 2.831180000000e-05, + 2.952830000000e-05, + 3.067910000000e-05, + 3.176630000000e-05, + 3.279220000000e-05,  \
+ 3.375920000000e-05, + 3.467000000000e-05, + 3.552700000000e-05, + 3.633260000000e-05, + 3.708950000000e-05,  \
+ 3.779990000000e-05, + 3.846610000000e-05, + 3.909060000000e-05, + 3.967550000000e-05, + 4.022310000000e-05,  \
+ 4.073550000000e-05, + 4.121500000000e-05, + 4.166370000000e-05, + 4.208360000000e-05, + 4.247670000000e-05,  \
+ 4.284510000000e-05, + 4.319060000000e-05, + 4.351490000000e-05, + 4.381970000000e-05, + 4.410660000000e-05,  \
+ 4.437690000000e-05, + 4.463200000000e-05, + 4.487330000000e-05, + 4.510170000000e-05, + 4.531830000000e-05,  \
+ 4.552420000000e-05, + 4.572010000000e-05, + 4.590690000000e-05, + 4.608520000000e-05, + 4.625580000000e-05,  \
+ 4.641930000000e-05, + 4.657610000000e-05, + 4.672680000000e-05, + 4.687190000000e-05, + 4.701170000000e-05,  \
+ 4.714670000000e-05, + 4.727710000000e-05, + 4.740330000000e-05, + 4.752560000000e-05, + 4.764430000000e-05,  \
+ 4.775950000000e-05, + 4.787160000000e-05, + 4.798060000000e-05, + 4.808680000000e-05, + 4.819040000000e-05,  \
+ 4.829160000000e-05, + 4.839040000000e-05, + 4.848700000000e-05, + 4.858150000000e-05, + 4.867410000000e-05,  \
+ 4.876490000000e-05, + 4.885390000000e-05, + 4.894120000000e-05, + 4.902700000000e-05, + 4.911130000000e-05,  \
+ 4.919410000000e-05, + 4.927570000000e-05, + 4.935590000000e-05, + 4.943490000000e-05, + 4.951280000000e-05 ]

.param id_pred_data_vg0.63=[ \
+ 2.189765073126e-06, + 4.331203526817e-06, + 6.422291044146e-06, + 8.461105171591e-06, + 1.044582822942e-05,  \
+ 1.237466902239e-05, + 1.424610061804e-05, + 1.605861471035e-05, + 1.781084094546e-05, + 1.950167352334e-05,  \
+ 2.113008042215e-05, + 2.269524615258e-05, + 2.419652315439e-05, + 2.563350659329e-05, + 2.700599652599e-05,  \
+ 2.831396181136e-05, + 2.955767384265e-05, + 3.073751810007e-05, + 3.185422639945e-05, + 3.290873137303e-05,  \
+ 3.390215453692e-05, + 3.483583423076e-05, + 3.571149703930e-05, + 3.653083811514e-05, + 3.729588206625e-05,  \
+ 3.800881240750e-05, + 3.867198349326e-05, + 3.928777063265e-05, + 3.985898889368e-05, + 4.038808256155e-05,  \
+ 4.087810579222e-05, + 4.133169073611e-05, + 4.175164227490e-05, + 4.214095592033e-05, + 4.250221099937e-05,  \
+ 4.283822810976e-05, + 4.315165126172e-05, + 4.344489527284e-05, + 4.372043105832e-05, + 4.398061428219e-05,  \
+ 4.422713580425e-05, + 4.446214545169e-05, + 4.468725805054e-05, + 4.490381776122e-05, + 4.511343286140e-05,  \
+ 4.531685815891e-05, + 4.551513426122e-05, + 4.570910241455e-05, + 4.589902455336e-05, + 4.608543895301e-05,  \
+ 4.626857349649e-05, + 4.644843807910e-05, + 4.662500723498e-05, + 4.679825957282e-05, + 4.696786854765e-05,  \
+ 4.713365691714e-05, + 4.729523090646e-05, + 4.745238780743e-05, + 4.760445066495e-05, + 4.775138804689e-05,  \
+ 4.789268787135e-05, + 4.802799987374e-05, + 4.815699554456e-05, + 4.827946890146e-05, + 4.839514331252e-05,  \
+ 4.850382407312e-05, + 4.860538458161e-05, + 4.869951779256e-05, + 4.878639374510e-05, + 4.886586757493e-05,  \
+ 4.893790268397e-05, + 4.900261759758e-05, + 4.906009686238e-05, + 4.911030919175e-05, + 4.915355930279e-05,  \
+ 4.918978753267e-05, + 4.921940337226e-05, + 4.924246619339e-05, + 4.925912828185e-05, + 4.926964757033e-05 ]

* Data table for Id-Vd at Vg = 0.64V
.param vd_data_vg0.64=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.64=[ \
+ 2.168900000000e-06, + 4.312600000000e-06, + 6.423700000000e-06, + 8.495300000000e-06, + 1.052110000000e-05,  \
+ 1.249570000000e-05, + 1.441420000000e-05, + 1.627260000000e-05, + 1.806780000000e-05, + 1.979730000000e-05,  \
+ 2.145930000000e-05, + 2.305250000000e-05, + 2.457620000000e-05, + 2.603040000000e-05, + 2.741530000000e-05,  \
+ 2.873180000000e-05, + 2.998120000000e-05, + 3.116500000000e-05, + 3.228520000000e-05, + 3.334400000000e-05,  \
+ 3.434350000000e-05, + 3.528640000000e-05, + 3.617510000000e-05, + 3.701190000000e-05, + 3.779940000000e-05,  \
+ 3.853980000000e-05, + 3.923550000000e-05, + 3.988880000000e-05, + 4.050170000000e-05, + 4.107660000000e-05,  \
+ 4.161550000000e-05, + 4.212050000000e-05, + 4.259370000000e-05, + 4.303720000000e-05, + 4.345300000000e-05,  \
+ 4.384290000000e-05, + 4.420880000000e-05, + 4.455250000000e-05, + 4.487570000000e-05, + 4.518000000000e-05,  \
+ 4.546670000000e-05, + 4.573730000000e-05, + 4.599310000000e-05, + 4.623530000000e-05, + 4.646490000000e-05,  \
+ 4.668290000000e-05, + 4.689030000000e-05, + 4.708790000000e-05, + 4.727650000000e-05, + 4.745670000000e-05,  \
+ 4.762920000000e-05, + 4.779460000000e-05, + 4.795340000000e-05, + 4.810610000000e-05, + 4.825320000000e-05,  \
+ 4.839500000000e-05, + 4.853200000000e-05, + 4.866440000000e-05, + 4.879260000000e-05, + 4.891680000000e-05,  \
+ 4.903740000000e-05, + 4.915450000000e-05, + 4.926840000000e-05, + 4.937930000000e-05, + 4.948730000000e-05,  \
+ 4.959270000000e-05, + 4.969550000000e-05, + 4.979600000000e-05, + 4.989430000000e-05, + 4.999050000000e-05,  \
+ 5.008470000000e-05, + 5.017700000000e-05, + 5.026750000000e-05, + 5.035630000000e-05, + 5.044360000000e-05,  \
+ 5.052930000000e-05, + 5.061360000000e-05, + 5.069650000000e-05, + 5.077810000000e-05, + 5.085840000000e-05 ]

.param id_pred_data_vg0.64=[ \
+ 2.207524812547e-06, + 4.367905203253e-06, + 6.479158764705e-06, + 8.539339760318e-06, + 1.054660824593e-05,  \
+ 1.249925378943e-05, + 1.439560655854e-05, + 1.623423187993e-05, + 1.801371050533e-05, + 1.973283360712e-05,  \
+ 2.139055446605e-05, + 2.298599516507e-05, + 2.451842694427e-05, + 2.598733728519e-05, + 2.739235424087e-05,  \
+ 2.873346908018e-05, + 3.001079952810e-05, + 3.122457215795e-05, + 3.237539771362e-05, + 3.346406447235e-05,  \
+ 3.449158000876e-05, + 3.545914136339e-05, + 3.636826048023e-05, + 3.722055698745e-05, + 3.801791535807e-05,  \
+ 3.876242466504e-05, + 3.945619959268e-05, + 4.010171629488e-05, + 4.070138369570e-05, + 4.125786654186e-05,  \
+ 4.177389622782e-05, + 4.225224256516e-05, + 4.269564058632e-05, + 4.310694523156e-05, + 4.348888032837e-05,  \
+ 4.384423722513e-05, + 4.417563621246e-05, + 4.448568128282e-05, + 4.477674207010e-05, + 4.505115794018e-05,  \
+ 4.531106962531e-05, + 4.555844425340e-05, + 4.579504522553e-05, + 4.602241358953e-05, + 4.624210523616e-05,  \
+ 4.645508903195e-05, + 4.666253254982e-05, + 4.686509608291e-05, + 4.706346080638e-05, + 4.725807593786e-05,  \
+ 4.744926365674e-05, + 4.763703153003e-05, + 4.782158466696e-05, + 4.800266833627e-05, + 4.818018278456e-05,  \
+ 4.835380124860e-05, + 4.852330741414e-05, + 4.868830699706e-05, + 4.884828951617e-05, + 4.900298954453e-05,  \
+ 4.915206962323e-05, + 4.929507587804e-05, + 4.943153136992e-05, + 4.956135991961e-05, + 4.968417633791e-05,  \
+ 4.979983787052e-05, + 4.990797024220e-05, + 5.000843870221e-05, + 5.010132968891e-05, + 5.018638912588e-05,  \
+ 5.026372826251e-05, + 5.033326568082e-05, + 5.039519332058e-05, + 5.044946417911e-05, + 5.049630090070e-05,  \
+ 5.053588363808e-05, + 5.056828063971e-05, + 5.059366871137e-05, + 5.061228373961e-05, + 5.062444251962e-05 ]

* Data table for Id-Vd at Vg = 0.65V
.param vd_data_vg0.65=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.65=[ \
+ 2.186800000000e-06, + 4.349200000000e-06, + 6.480000000000e-06, + 8.572200000000e-06, + 1.061980000000e-05,  \
+ 1.261720000000e-05, + 1.455950000000e-05, + 1.644300000000e-05, + 1.826420000000e-05, + 2.002080000000e-05,  \
+ 2.171080000000e-05, + 2.333290000000e-05, + 2.488640000000e-05, + 2.637100000000e-05, + 2.778700000000e-05,  \
+ 2.913510000000e-05, + 3.041630000000e-05, + 3.163220000000e-05, + 3.278440000000e-05, + 3.387500000000e-05,  \
+ 3.490620000000e-05, + 3.588050000000e-05, + 3.680000000000e-05, + 3.766730000000e-05, + 3.848480000000e-05,  \
+ 3.925470000000e-05, + 3.997930000000e-05, + 4.066080000000e-05, + 4.130140000000e-05, + 4.190320000000e-05,  \
+ 4.246830000000e-05, + 4.299870000000e-05, + 4.349650000000e-05, + 4.396360000000e-05, + 4.440200000000e-05,  \
+ 4.481360000000e-05, + 4.520030000000e-05, + 4.556370000000e-05, + 4.590560000000e-05, + 4.622760000000e-05,  \
+ 4.653120000000e-05, + 4.681770000000e-05, + 4.708850000000e-05, + 4.734480000000e-05, + 4.758770000000e-05,  \
+ 4.781840000000e-05, + 4.803760000000e-05, + 4.824640000000e-05, + 4.844550000000e-05, + 4.863570000000e-05,  \
+ 4.881760000000e-05, + 4.899190000000e-05, + 4.915920000000e-05, + 4.931980000000e-05, + 4.947450000000e-05,  \
+ 4.962340000000e-05, + 4.976710000000e-05, + 4.990600000000e-05, + 5.004030000000e-05, + 5.017030000000e-05,  \
+ 5.029640000000e-05, + 5.041880000000e-05, + 5.053780000000e-05, + 5.065340000000e-05, + 5.076600000000e-05,  \
+ 5.087580000000e-05, + 5.098290000000e-05, + 5.108740000000e-05, + 5.118950000000e-05, + 5.128940000000e-05,  \
+ 5.138710000000e-05, + 5.148280000000e-05, + 5.157670000000e-05, + 5.166870000000e-05, + 5.175900000000e-05,  \
+ 5.184760000000e-05, + 5.193470000000e-05, + 5.202040000000e-05, + 5.210460000000e-05, + 5.218750000000e-05 ]

.param id_pred_data_vg0.65=[ \
+ 2.224314666819e-06, + 4.402603954077e-06, + 6.532890693052e-06, + 8.613269310445e-06, + 1.064189273166e-05,  \
+ 1.261705270736e-05, + 1.453708566260e-05, + 1.640047412366e-05, + 1.820584599045e-05, + 1.995192287723e-05,  \
+ 2.163762255805e-05, + 2.326196059585e-05, + 2.482419789885e-05, + 2.632372692460e-05, + 2.776011024253e-05,  \
+ 2.913320204243e-05, + 3.044296201551e-05, + 3.168968134560e-05, + 3.287366489531e-05, + 3.399558481760e-05,  \
+ 3.505640241201e-05, + 3.605720208725e-05, + 3.699925917317e-05, + 3.788404050283e-05, + 3.871340595651e-05,  \
+ 3.948911733460e-05, + 4.021341941552e-05, + 4.088848072570e-05, + 4.151673638262e-05, + 4.210070183035e-05,  \
+ 4.264304865501e-05, + 4.314632620662e-05, + 4.361345287180e-05, + 4.404712264659e-05, + 4.445015001693e-05,  \
+ 4.482528136577e-05, + 4.517503955867e-05, + 4.550220837700e-05, + 4.580918015563e-05, + 4.609840980265e-05,  \
+ 4.637196761905e-05, + 4.663207131671e-05, + 4.688037173764e-05, + 4.711883637356e-05, + 4.734877184092e-05,  \
+ 4.757143760798e-05, + 4.778805501701e-05, + 4.799939808436e-05, + 4.820628826565e-05, + 4.840908877668e-05,  \
+ 4.860827197263e-05, + 4.880407417659e-05, + 4.899650921288e-05, + 4.918546750559e-05, + 4.937083940604e-05,  \
+ 4.955238720868e-05, + 4.972979309969e-05, + 4.990270390408e-05, + 5.007068575651e-05, + 5.023337871535e-05,  \
+ 5.039028495958e-05, + 5.054113920778e-05, + 5.068543985544e-05, + 5.082292016596e-05, + 5.095319465909e-05,  \
+ 5.107589400723e-05, + 5.119119283336e-05, + 5.129840516020e-05, + 5.139761480677e-05, + 5.148874843144e-05,  \
+ 5.157183470146e-05, + 5.164667847566e-05, + 5.171352684556e-05, + 5.177237500902e-05, + 5.182326094655e-05,  \
+ 5.186645226786e-05, + 5.190213203605e-05, + 5.193036529818e-05, + 5.195146004553e-05, + 5.196561687626e-05 ]

* Data table for Id-Vd at Vg = 0.66V
.param vd_data_vg0.66=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.66=[ \
+ 2.204000000000e-06, + 4.384300000000e-06, + 6.533900000000e-06, + 8.646000000000e-06, + 1.071440000000e-05,  \
+ 1.273360000000e-05, + 1.469880000000e-05, + 1.660620000000e-05, + 1.845240000000e-05, + 2.023500000000e-05,  \
+ 2.195190000000e-05, + 2.360180000000e-05, + 2.518390000000e-05, + 2.669790000000e-05, + 2.814380000000e-05,  \
+ 2.952230000000e-05, + 3.083430000000e-05, + 3.208110000000e-05, + 3.326430000000e-05, + 3.438590000000e-05,  \
+ 3.544790000000e-05, + 3.645260000000e-05, + 3.740240000000e-05, + 3.829940000000e-05, + 3.914620000000e-05,  \
+ 3.994490000000e-05, + 4.069780000000e-05, + 4.140710000000e-05, + 4.207480000000e-05, + 4.270320000000e-05,  \
+ 4.329410000000e-05, + 4.384970000000e-05, + 4.437190000000e-05, + 4.486250000000e-05, + 4.532360000000e-05,  \
+ 4.575700000000e-05, + 4.616450000000e-05, + 4.654790000000e-05, + 4.690880000000e-05, + 4.724880000000e-05,  \
+ 4.756950000000e-05, + 4.787220000000e-05, + 4.815840000000e-05, + 4.842920000000e-05, + 4.868590000000e-05,  \
+ 4.892950000000e-05, + 4.916100000000e-05, + 4.938130000000e-05, + 4.959140000000e-05, + 4.979180000000e-05,  \
+ 4.998350000000e-05, + 5.016700000000e-05, + 5.034300000000e-05, + 5.051190000000e-05, + 5.067430000000e-05,  \
+ 5.083070000000e-05, + 5.098140000000e-05, + 5.112690000000e-05, + 5.126760000000e-05, + 5.140370000000e-05,  \
+ 5.153550000000e-05, + 5.166340000000e-05, + 5.178750000000e-05, + 5.190810000000e-05, + 5.202550000000e-05,  \
+ 5.213980000000e-05, + 5.225120000000e-05, + 5.235990000000e-05, + 5.246600000000e-05, + 5.256970000000e-05,  \
+ 5.267110000000e-05, + 5.277040000000e-05, + 5.286760000000e-05, + 5.296280000000e-05, + 5.305630000000e-05,  \
+ 5.314800000000e-05, + 5.323800000000e-05, + 5.332650000000e-05, + 5.341340000000e-05, + 5.349890000000e-05 ]

.param id_pred_data_vg0.66=[ \
+ 2.240150934085e-06, + 4.435340233613e-06, + 6.583595095435e-06, + 8.683026535437e-06, + 1.073182502296e-05,  \
+ 1.272827532375e-05, + 1.467068970669e-05, + 1.655759755522e-05, + 1.838754207711e-05, + 2.015925274463e-05,  \
+ 2.187160323956e-05, + 2.352353185415e-05, + 2.511432598112e-05, + 2.664319297764e-05, + 2.810971418512e-05,  \
+ 2.951360540465e-05, + 3.085470554652e-05, + 3.213320713257e-05, + 3.334937355248e-05, + 3.450371441431e-05,  \
+ 3.559704957297e-05, + 3.663025971036e-05, + 3.760460691410e-05, + 3.852142137475e-05, + 3.938231020584e-05,  \
+ 4.018901527161e-05, + 4.094360760064e-05, + 4.164815763943e-05, + 4.230490347254e-05, + 4.291649238439e-05,  \
+ 4.348510294221e-05, + 4.401372279972e-05, + 4.450483422261e-05, + 4.496117646340e-05, + 4.538567372947e-05,  \
+ 4.578079737257e-05, + 4.614940902684e-05, + 4.649413924199e-05, + 4.681744736445e-05, + 4.712171503343e-05,  \
+ 4.740939126350e-05, + 4.768245518790e-05, + 4.794288404810e-05, + 4.819254507311e-05, + 4.843294154853e-05,  \
+ 4.866548551945e-05, + 4.889137337159e-05, + 4.911162424833e-05, + 4.932697571348e-05, + 4.953808092978e-05,  \
+ 4.974523108103e-05, + 4.994894552510e-05, + 5.014924485295e-05, + 5.034610701841e-05, + 5.053927416157e-05,  \
+ 5.072864878457e-05, + 5.091405342682e-05, + 5.109492863994e-05, + 5.127093536430e-05, + 5.144164751982e-05,  \
+ 5.160661043192e-05, + 5.176549966563e-05, + 5.191780423047e-05, + 5.206304602325e-05, + 5.220102539170e-05,  \
+ 5.233147385297e-05, + 5.245390675555e-05, + 5.256817530608e-05, + 5.267426007777e-05, + 5.277188611217e-05,  \
+ 5.286102867103e-05, + 5.294178205077e-05, + 5.301389173837e-05, + 5.307771178195e-05, + 5.313327710610e-05,  \
+ 5.318055336829e-05, + 5.321992670360e-05, + 5.325146630639e-05, + 5.327548460627e-05, + 5.329204141162e-05 ]

* Data table for Id-Vd at Vg = 0.67V
.param vd_data_vg0.67=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.67=[ \
+ 2.220400000000e-06, + 4.418000000000e-06, + 6.585600000000e-06, + 8.716700000000e-06, + 1.080500000000e-05,  \
+ 1.284510000000e-05, + 1.483240000000e-05, + 1.676270000000e-05, + 1.863290000000e-05, + 2.044030000000e-05,  \
+ 2.218300000000e-05, + 2.385970000000e-05, + 2.546920000000e-05, + 2.701140000000e-05, + 2.848620000000e-05,  \
+ 2.989390000000e-05, + 3.123560000000e-05, + 3.251230000000e-05, + 3.372560000000e-05, + 3.487720000000e-05,  \
+ 3.596920000000e-05, + 3.700360000000e-05, + 3.798260000000e-05, + 3.890870000000e-05, + 3.978400000000e-05,  \
+ 4.061090000000e-05, + 4.139140000000e-05, + 4.212790000000e-05, + 4.282230000000e-05, + 4.347670000000e-05,  \
+ 4.409320000000e-05, + 4.467360000000e-05, + 4.521990000000e-05, + 4.573390000000e-05, + 4.621760000000e-05,  \
+ 4.667280000000e-05, + 4.710120000000e-05, + 4.750460000000e-05, + 4.788470000000e-05, + 4.824290000000e-05,  \
+ 4.858100000000e-05, + 4.890020000000e-05, + 4.920210000000e-05, + 4.948770000000e-05, + 4.975850000000e-05,  \
+ 5.001540000000e-05, + 5.025940000000e-05, + 5.049170000000e-05, + 5.071300000000e-05, + 5.092410000000e-05,  \
+ 5.112580000000e-05, + 5.131880000000e-05, + 5.150380000000e-05, + 5.168120000000e-05, + 5.185170000000e-05,  \
+ 5.201580000000e-05, + 5.217380000000e-05, + 5.232620000000e-05, + 5.247340000000e-05, + 5.261570000000e-05,  \
+ 5.275350000000e-05, + 5.288700000000e-05, + 5.301650000000e-05, + 5.314230000000e-05, + 5.326460000000e-05,  \
+ 5.338360000000e-05, + 5.349950000000e-05, + 5.361240000000e-05, + 5.372270000000e-05, + 5.383030000000e-05,  \
+ 5.393550000000e-05, + 5.403840000000e-05, + 5.413910000000e-05, + 5.423770000000e-05, + 5.433440000000e-05,  \
+ 5.442920000000e-05, + 5.452220000000e-05, + 5.461360000000e-05, + 5.470340000000e-05, + 5.479160000000e-05 ]

.param id_pred_data_vg0.67=[ \
+ 2.255063009216e-06, + 4.466147220228e-06, + 6.631333963014e-06, + 8.748741820455e-06, + 1.081657319446e-05,  \
+ 1.283310935833e-05, + 1.479671409470e-05, + 1.670588389970e-05, + 1.855911832536e-05, + 2.035520155914e-05,  \
+ 2.209291749750e-05, + 2.377119439188e-05, + 2.538921980886e-05, + 2.694622846320e-05, + 2.844165937859e-05,  \
+ 2.987511688843e-05, + 3.124649767415e-05, + 3.255569958128e-05, + 3.380306836334e-05, + 3.498892474454e-05,  \
+ 3.611389125581e-05, + 3.717879764736e-05, + 3.818477227469e-05, + 3.913300693966e-05, + 4.002493005828e-05,  \
+ 4.086233035196e-05, + 4.164687808952e-05, + 4.238070629071e-05, + 4.306596092647e-05, + 4.370505484985e-05,  \
+ 4.430020795553e-05, + 4.485417157412e-05, + 4.536950131296e-05, + 4.584891867125e-05, + 4.629508475773e-05,  \
+ 4.671068571042e-05, + 4.709846194601e-05, + 4.746105085360e-05, + 4.780106697581e-05, + 4.812085826416e-05,  \
+ 4.842289905355e-05, + 4.870927805314e-05, + 4.898209095700e-05, + 4.924317472614e-05, + 4.949423782818e-05,  \
+ 4.973680770490e-05, + 4.997210460715e-05, + 5.020129261538e-05, + 5.042517019319e-05, + 5.064440847491e-05,  \
+ 5.085986638733e-05, + 5.107141099870e-05, + 5.127948694280e-05, + 5.148402502527e-05, + 5.168495881662e-05,  \
+ 5.188228853513e-05, + 5.207553680521e-05, + 5.226432709605e-05, + 5.244836436759e-05, + 5.262721097097e-05,  \
+ 5.280035809847e-05, + 5.296726405504e-05, + 5.312761146342e-05, + 5.328101571649e-05, + 5.342696385924e-05,  \
+ 5.356517518521e-05, + 5.369530765165e-05, + 5.381699709687e-05, + 5.393023129727e-05, + 5.403477844084e-05,  \
+ 5.413048878836e-05, + 5.421736626886e-05, + 5.429541160993e-05, + 5.436461302452e-05, + 5.442520341603e-05,  \
+ 5.447716946946e-05, + 5.452072342450e-05, + 5.455600126879e-05, + 5.458331128466e-05, + 5.460293032229e-05 ]

* Data table for Id-Vd at Vg = 0.68V
.param vd_data_vg0.68=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.68=[ \
+ 2.236200000000e-06, + 4.450300000000e-06, + 6.635200000000e-06, + 8.784500000000e-06, + 1.089190000000e-05,  \
+ 1.295210000000e-05, + 1.496040000000e-05, + 1.691270000000e-05, + 1.880590000000e-05, + 2.063720000000e-05,  \
+ 2.240470000000e-05, + 2.410700000000e-05, + 2.574300000000e-05, + 2.731220000000e-05, + 2.881470000000e-05,  \
+ 3.025070000000e-05, + 3.162100000000e-05, + 3.292660000000e-05, + 3.416890000000e-05, + 3.534960000000e-05,  \
+ 3.647060000000e-05, + 3.753380000000e-05, + 3.854140000000e-05, + 3.949570000000e-05, + 4.039890000000e-05,  \
+ 4.125310000000e-05, + 4.206070000000e-05, + 4.282370000000e-05, + 4.354420000000e-05, + 4.422420000000e-05,  \
+ 4.486570000000e-05, + 4.547050000000e-05, + 4.604060000000e-05, + 4.657780000000e-05, + 4.708390000000e-05,  \
+ 4.756080000000e-05, + 4.801010000000e-05, + 4.843360000000e-05, + 4.883280000000e-05, + 4.920950000000e-05,  \
+ 4.956510000000e-05, + 4.990110000000e-05, + 5.021890000000e-05, + 5.051970000000e-05, + 5.080470000000e-05,  \
+ 5.107520000000e-05, + 5.133220000000e-05, + 5.157660000000e-05, + 5.180940000000e-05, + 5.203150000000e-05,  \
+ 5.224350000000e-05, + 5.244640000000e-05, + 5.264060000000e-05, + 5.282680000000e-05, + 5.300570000000e-05,  \
+ 5.317760000000e-05, + 5.334310000000e-05, + 5.350270000000e-05, + 5.365660000000e-05, + 5.380540000000e-05,  \
+ 5.394930000000e-05, + 5.408860000000e-05, + 5.422370000000e-05, + 5.435480000000e-05, + 5.448220000000e-05,  \
+ 5.460600000000e-05, + 5.472650000000e-05, + 5.484390000000e-05, + 5.495840000000e-05, + 5.507010000000e-05,  \
+ 5.517920000000e-05, + 5.528590000000e-05, + 5.539020000000e-05, + 5.549230000000e-05, + 5.559230000000e-05,  \
+ 5.569030000000e-05, + 5.578640000000e-05, + 5.588070000000e-05, + 5.597340000000e-05, + 5.606440000000e-05 ]

.param id_pred_data_vg0.68=[ \
+ 2.269070246257e-06, + 4.495097091421e-06, + 6.676190241706e-06, + 8.810517028905e-06, + 1.089627403417e-05,  \
+ 1.293176261242e-05, + 1.491536866524e-05, + 1.684556598775e-05, + 1.872091917903e-05, + 2.054010401480e-05,  \
+ 2.230191908893e-05, + 2.400531840976e-05, + 2.564933151007e-05, + 2.723322249949e-05, + 2.875634309021e-05,  \
+ 3.021828364581e-05, + 3.161877131788e-05, + 3.295767994132e-05, + 3.423517235206e-05, + 3.545157087501e-05,  \
+ 3.660729111289e-05, + 3.770317445742e-05, + 3.874003639794e-05, + 3.971909754910e-05, + 4.064158565598e-05,  \
+ 4.150918364758e-05, + 4.232346269418e-05, + 4.308634262998e-05, + 4.379996360512e-05, + 4.446644161362e-05,  \
+ 4.508821482887e-05, + 4.566770978272e-05, + 4.620749736205e-05, + 4.671002272516e-05, + 4.717824558611e-05,  \
+ 4.761457967106e-05, + 4.802189680049e-05, + 4.840281879297e-05, + 4.875980346696e-05, + 4.909542039968e-05,  \
+ 4.941215687722e-05, + 4.971220681909e-05, + 4.999769211281e-05, + 5.027046921896e-05, + 5.053240856796e-05,  \
+ 5.078520000097e-05, + 5.103002986289e-05, + 5.126817617565e-05, + 5.150069344381e-05, + 5.172830788069e-05,  \
+ 5.195154706598e-05, + 5.217096739216e-05, + 5.238672260020e-05, + 5.259908793960e-05, + 5.280774530547e-05,  \
+ 5.301280121785e-05, + 5.321380776877e-05, + 5.341059542843e-05, + 5.360265509808e-05, + 5.378959758673e-05,  \
+ 5.397084001743e-05, + 5.414599028882e-05, + 5.431461861008e-05, + 5.447617731988e-05, + 5.463024390338e-05,  \
+ 5.477647937369e-05, + 5.491447904205e-05, + 5.504397006007e-05, + 5.516468001588e-05, + 5.527641187655e-05,  \
+ 5.537907338294e-05, + 5.547266628128e-05, + 5.555697105592e-05, + 5.563213111600e-05, + 5.569817221840e-05,  \
+ 5.575522780418e-05, + 5.580337368883e-05, + 5.584304512013e-05, + 5.587409512373e-05, + 5.589705542661e-05 ]

* Data table for Id-Vd at Vg = 0.69V
.param vd_data_vg0.69=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.69=[ \
+ 2.251400000000e-06, + 4.481200000000e-06, + 6.682800000000e-06, + 8.849500000000e-06, + 1.097520000000e-05,  \
+ 1.305470000000e-05, + 1.508310000000e-05, + 1.705660000000e-05, + 1.897180000000e-05, + 2.082610000000e-05,  \
+ 2.261740000000e-05, + 2.434420000000e-05, + 2.600560000000e-05, + 2.760090000000e-05, + 2.913000000000e-05,  \
+ 3.059320000000e-05, + 3.199100000000e-05, + 3.332450000000e-05, + 3.459490000000e-05, + 3.580370000000e-05,  \
+ 3.695270000000e-05, + 3.804390000000e-05, + 3.907920000000e-05, + 4.006100000000e-05, + 4.099120000000e-05,  \
+ 4.187230000000e-05, + 4.270620000000e-05, + 4.349510000000e-05, + 4.424100000000e-05, + 4.494600000000e-05,  \
+ 4.561190000000e-05, + 4.624070000000e-05, + 4.683420000000e-05, + 4.739420000000e-05, + 4.792260000000e-05,  \
+ 4.842090000000e-05, + 4.889100000000e-05, + 4.933450000000e-05, + 4.975300000000e-05, + 5.014820000000e-05,  \
+ 5.052150000000e-05, + 5.087440000000e-05, + 5.120820000000e-05, + 5.152430000000e-05, + 5.182400000000e-05,  \
+ 5.210830000000e-05, + 5.237840000000e-05, + 5.263530000000e-05, + 5.287990000000e-05, + 5.311320000000e-05,  \
+ 5.333590000000e-05, + 5.354870000000e-05, + 5.375250000000e-05, + 5.394780000000e-05, + 5.413520000000e-05,  \
+ 5.431530000000e-05, + 5.448850000000e-05, + 5.465540000000e-05, + 5.481630000000e-05, + 5.497170000000e-05,  \
+ 5.512200000000e-05, + 5.526730000000e-05, + 5.540810000000e-05, + 5.554470000000e-05, + 5.567730000000e-05,  \
+ 5.580610000000e-05, + 5.593140000000e-05, + 5.605340000000e-05, + 5.617220000000e-05, + 5.628820000000e-05,  \
+ 5.640130000000e-05, + 5.651180000000e-05, + 5.661980000000e-05, + 5.672540000000e-05, + 5.682880000000e-05,  \
+ 5.693010000000e-05, + 5.702940000000e-05, + 5.712680000000e-05, + 5.722240000000e-05, + 5.731620000000e-05 ]

.param id_pred_data_vg0.69=[ \
+ 2.282193454448e-06, + 4.522241652012e-06, + 6.718261283822e-06, + 8.868464501575e-06, + 1.097108906833e-05,  \
+ 1.302444026805e-05, + 1.502690502093e-05, + 1.697700703517e-05, + 1.887325634016e-05, + 2.071433409583e-05,  \
+ 2.249903220218e-05, + 2.422628807835e-05, + 2.589508862002e-05, + 2.750467217993e-05, + 2.905433284468e-05,  \
+ 3.054356435314e-05, + 3.197205587639e-05, + 3.333955944981e-05, + 3.464619425358e-05, + 3.589218249545e-05,  \
+ 3.707785726874e-05, + 3.820374869974e-05, + 3.927084777388e-05, + 4.028007388115e-05, + 4.123265171074e-05,  \
+ 4.212993837427e-05, + 4.297352250433e-05, + 4.376527038403e-05, + 4.450702967006e-05, + 4.520098445937e-05,  \
+ 4.584915965097e-05, + 4.645424894989e-05, + 4.701849102275e-05, + 4.754452325869e-05, + 4.803494230146e-05,  \
+ 4.849242162891e-05, + 4.891951975878e-05, + 4.931903386023e-05, + 4.969344401616e-05, + 5.004536360502e-05,  \
+ 5.037711103796e-05, + 5.069104896393e-05, + 5.098939967866e-05, + 5.127418844495e-05, + 5.154740138096e-05,  \
+ 5.181041473406e-05, + 5.206495079619e-05, + 5.231221555732e-05, + 5.255327807390e-05, + 5.278916796669e-05,  \
+ 5.302047720761e-05, + 5.324766010744e-05, + 5.347102895030e-05, + 5.369091071771e-05, + 5.390729747887e-05,  \
+ 5.411997495685e-05, + 5.432870457298e-05, + 5.453330741148e-05, + 5.473326666106e-05, + 5.492828786373e-05,  \
+ 5.511767893040e-05, + 5.530113703571e-05, + 5.547796848987e-05, + 5.564792081714e-05, + 5.581025070569e-05,  \
+ 5.596471411991e-05, + 5.611084568955e-05, + 5.624836194329e-05, + 5.637681802909e-05, + 5.649623126374e-05,  \
+ 5.660623486619e-05, + 5.670677055605e-05, + 5.679771493305e-05, + 5.687916229363e-05, + 5.695124491467e-05,  \
+ 5.701383255655e-05, + 5.706714357075e-05, + 5.711147416150e-05, + 5.714698541851e-05, + 5.717368912883e-05 ]

* Data table for Id-Vd at Vg = 0.70V
.param vd_data_vg0.70=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.70=[ \
+ 2.265900000000e-06, + 4.511000000000e-06, + 6.728400000000e-06, + 8.911800000000e-06, + 1.105520000000e-05,  \
+ 1.315310000000e-05, + 1.520090000000e-05, + 1.719470000000e-05, + 1.913100000000e-05, + 2.100730000000e-05,  \
+ 2.282140000000e-05, + 2.457190000000e-05, + 2.625760000000e-05, + 2.787790000000e-05, + 2.943260000000e-05,  \
+ 3.092190000000e-05, + 3.234630000000e-05, + 3.370660000000e-05, + 3.500410000000e-05, + 3.624010000000e-05,  \
+ 3.741630000000e-05, + 3.853450000000e-05, + 3.959680000000e-05, + 4.060510000000e-05, + 4.156170000000e-05,  \
+ 4.246870000000e-05, + 4.332820000000e-05, + 4.414240000000e-05, + 4.491310000000e-05, + 4.564250000000e-05,  \
+ 4.633240000000e-05, + 4.698460000000e-05, + 4.760110000000e-05, + 4.818350000000e-05, + 4.873370000000e-05,  \
+ 4.925320000000e-05, + 4.974390000000e-05, + 5.020730000000e-05, + 5.064510000000e-05, + 5.105870000000e-05,  \
+ 5.144970000000e-05, + 5.181950000000e-05, + 5.216960000000e-05, + 5.250120000000e-05, + 5.281560000000e-05,  \
+ 5.311400000000e-05, + 5.339740000000e-05, + 5.366700000000e-05, + 5.392370000000e-05, + 5.416840000000e-05,  \
+ 5.440190000000e-05, + 5.462510000000e-05, + 5.483860000000e-05, + 5.504320000000e-05, + 5.523940000000e-05,  \
+ 5.542780000000e-05, + 5.560900000000e-05, + 5.578350000000e-05, + 5.595160000000e-05, + 5.611380000000e-05,  \
+ 5.627050000000e-05, + 5.642210000000e-05, + 5.656880000000e-05, + 5.671100000000e-05, + 5.684890000000e-05,  \
+ 5.698290000000e-05, + 5.711310000000e-05, + 5.723980000000e-05, + 5.736310000000e-05, + 5.748330000000e-05,  \
+ 5.760060000000e-05, + 5.771500000000e-05, + 5.782680000000e-05, + 5.793610000000e-05, + 5.804310000000e-05,  \
+ 5.814780000000e-05, + 5.825030000000e-05, + 5.835080000000e-05, + 5.844940000000e-05, + 5.854620000000e-05 ]

.param id_pred_data_vg0.70=[ \
+ 2.294464648003e-06, + 4.547615535557e-06, + 6.757625669707e-06, + 8.922707638703e-06, + 1.104117181967e-05,  \
+ 1.311130385147e-05, + 1.513155235443e-05, + 1.710038864985e-05, + 1.901640091091e-05, + 2.087821194436e-05,  \
+ 2.268468582770e-05, + 2.443458361086e-05, + 2.612704920466e-05, + 2.776110923151e-05, + 2.933612631750e-05,  \
+ 3.085151081905e-05, + 3.230691043427e-05, + 3.370200865902e-05, + 3.503677828121e-05, + 3.631132130977e-05,  \
+ 3.752601143788e-05, + 3.868125990266e-05, + 3.977774191299e-05, + 4.081653314643e-05, + 4.179845564067e-05,  \
+ 4.272496153135e-05, + 4.359750542790e-05, + 4.441768920515e-05, + 4.518734902376e-05, + 4.590850876411e-05,  \
+ 4.658321835450e-05, + 4.721384029835e-05, + 4.780275601661e-05, + 4.835236584768e-05, + 4.886519018328e-05,  \
+ 4.934403346851e-05, + 4.979130928405e-05, + 5.020967393648e-05, + 5.060189214419e-05, + 5.097026005387e-05,  \
+ 5.131739162607e-05, + 5.164560279809e-05, + 5.195720739721e-05, + 5.225432600128e-05, + 5.253872514004e-05,  \
+ 5.281233476126e-05, + 5.307665196597e-05, + 5.333314882591e-05, + 5.358295260521e-05, + 5.382710878621e-05,  \
+ 5.406626347394e-05, + 5.430119024822e-05, + 5.453225559904e-05, + 5.475958372699e-05, + 5.498336722667e-05,  \
+ 5.520355713088e-05, + 5.542000326386e-05, + 5.563227314269e-05, + 5.584015183558e-05, + 5.604306788882e-05,  \
+ 5.624064848234e-05, + 5.643225769745e-05, + 5.661740440701e-05, + 5.679566878825e-05, + 5.696639782400e-05,  \
+ 5.712923593819e-05, + 5.728375923354e-05, + 5.742946523242e-05, + 5.756605292845e-05, + 5.769332492491e-05,  \
+ 5.781095038401e-05, + 5.791881470941e-05, + 5.801690494991e-05, + 5.810519505758e-05, + 5.818360841658e-05,  \
+ 5.825220956467e-05, + 5.831118709466e-05, + 5.836060168804e-05, + 5.840084406373e-05, + 5.843203398399e-05 ]

* Data table for Id-Vd at Vg = 0.71V
.param vd_data_vg0.71=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.71=[ \
+ 2.279900000000e-06, + 4.539500000000e-06, + 6.772300000000e-06, + 8.971700000000e-06, + 1.113190000000e-05,  \
+ 1.324760000000e-05, + 1.531400000000e-05, + 1.732710000000e-05, + 1.928380000000e-05, + 2.118120000000e-05,  \
+ 2.301720000000e-05, + 2.479030000000e-05, + 2.649940000000e-05, + 2.814370000000e-05, + 2.972300000000e-05,  \
+ 3.123740000000e-05, + 3.268730000000e-05, + 3.407350000000e-05, + 3.539710000000e-05, + 3.665930000000e-05,  \
+ 3.786180000000e-05, + 3.900620000000e-05, + 4.009450000000e-05, + 4.112870000000e-05, + 4.211090000000e-05,  \
+ 4.304310000000e-05, + 4.392750000000e-05, + 4.476620000000e-05, + 4.556110000000e-05, + 4.631420000000e-05,  \
+ 4.702740000000e-05, + 4.770250000000e-05, + 4.834150000000e-05, + 4.894590000000e-05, + 4.951750000000e-05,  \
+ 5.005790000000e-05, + 5.056890000000e-05, + 5.105200000000e-05, + 5.150880000000e-05, + 5.194080000000e-05,  \
+ 5.234950000000e-05, + 5.273640000000e-05, + 5.310270000000e-05, + 5.344990000000e-05, + 5.377920000000e-05,  \
+ 5.409170000000e-05, + 5.438870000000e-05, + 5.467120000000e-05, + 5.494010000000e-05, + 5.519640000000e-05,  \
+ 5.544100000000e-05, + 5.567470000000e-05, + 5.589820000000e-05, + 5.611230000000e-05, + 5.631750000000e-05,  \
+ 5.651450000000e-05, + 5.670380000000e-05, + 5.688600000000e-05, + 5.706140000000e-05, + 5.723070000000e-05,  \
+ 5.739400000000e-05, + 5.755200000000e-05, + 5.770470000000e-05, + 5.785270000000e-05, + 5.799620000000e-05,  \
+ 5.813540000000e-05, + 5.827070000000e-05, + 5.840220000000e-05, + 5.853010000000e-05, + 5.865480000000e-05,  \
+ 5.877620000000e-05, + 5.889480000000e-05, + 5.901050000000e-05, + 5.912350000000e-05, + 5.923400000000e-05,  \
+ 5.934220000000e-05, + 5.944800000000e-05, + 5.955180000000e-05, + 5.965340000000e-05, + 5.975320000000e-05 ]

.param id_pred_data_vg0.71=[ \
+ 2.305899979547e-06, + 4.571282770485e-06, + 6.794355867896e-06, + 8.973396616057e-06, + 1.110668090405e-05,  \
+ 1.319259259617e-05, + 1.522954902612e-05, + 1.721607754007e-05, + 1.915071305120e-05, + 2.103213191731e-05,  \
+ 2.285918089910e-05, + 2.463061886374e-05, + 2.634552918607e-05, + 2.800302667310e-05, + 2.960224301205e-05,  \
+ 3.114268649369e-05, + 3.262385944254e-05, + 3.404546761885e-05, + 3.540734469425e-05, + 3.670950827654e-05,  \
+ 3.795228229137e-05, + 3.913595457561e-05, + 4.026114052976e-05, + 4.132867092267e-05, + 4.233951040078e-05,  \
+ 4.329468443757e-05, + 4.419563541887e-05, + 4.504394950345e-05, + 4.584124661051e-05, + 4.658949910663e-05,  \
+ 4.729049469461e-05, + 4.794664680958e-05, + 4.856031155214e-05, + 4.913352575386e-05, + 4.966908090864e-05,  \
+ 5.016938899644e-05, + 5.063708769740e-05, + 5.107468372444e-05, + 5.148490381544e-05, + 5.187008646317e-05,  \
+ 5.223295986070e-05, + 5.257584998617e-05, + 5.290088374750e-05, + 5.321045609890e-05, + 5.350648789317e-05,  \
+ 5.379077600082e-05, + 5.406520176621e-05, + 5.433098296635e-05, + 5.458951738547e-05, + 5.484186840476e-05,  \
+ 5.508905429451e-05, + 5.533174698940e-05, + 5.557016731473e-05, + 5.580496159382e-05, + 5.603611862171e-05,  \
+ 5.626369034871e-05, + 5.648757942254e-05, + 5.670745464158e-05, + 5.692303588148e-05, + 5.713381542591e-05,  \
+ 5.733939360653e-05, + 5.753913574154e-05, + 5.773259174020e-05, + 5.791928619146e-05, + 5.809849135403e-05,  \
+ 5.826979031553e-05, + 5.843274680956e-05, + 5.858690390596e-05, + 5.873179230548e-05, + 5.886719882255e-05,  \
+ 5.899278599827e-05, + 5.910849489737e-05, + 5.921390373260e-05, + 5.930933562922e-05, + 5.939458606008e-05,  \
+ 5.946960678557e-05, + 5.953458545264e-05, + 5.958969559288e-05, + 5.963516523479e-05, + 5.967110628262e-05 ]

* Data table for Id-Vd at Vg = 0.72V
.param vd_data_vg0.72=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.72=[ \
+ 2.293300000000e-06, + 4.566900000000e-06, + 6.814400000000e-06, + 9.029200000000e-06, + 1.120560000000e-05,  \
+ 1.333830000000e-05, + 1.542250000000e-05, + 1.745430000000e-05, + 1.943040000000e-05, + 2.134810000000e-05,  \
+ 2.320510000000e-05, + 2.500000000000e-05, + 2.673150000000e-05, + 2.839880000000e-05, + 3.000180000000e-05,  \
+ 3.154030000000e-05, + 3.301480000000e-05, + 3.442590000000e-05, + 3.577450000000e-05, + 3.706200000000e-05,  \
+ 3.828980000000e-05, + 3.945960000000e-05, + 4.057310000000e-05, + 4.163230000000e-05, + 4.263930000000e-05,  \
+ 4.359600000000e-05, + 4.450460000000e-05, + 4.536700000000e-05, + 4.618540000000e-05, + 4.696160000000e-05,  \
+ 4.769750000000e-05, + 4.839490000000e-05, + 4.905580000000e-05, + 4.968160000000e-05, + 5.027420000000e-05,  \
+ 5.083520000000e-05, + 5.136610000000e-05, + 5.186870000000e-05, + 5.234430000000e-05, + 5.279450000000e-05,  \
+ 5.322080000000e-05, + 5.362460000000e-05, + 5.400720000000e-05, + 5.437000000000e-05, + 5.471420000000e-05,  \
+ 5.504110000000e-05, + 5.535170000000e-05, + 5.564720000000e-05, + 5.592850000000e-05, + 5.619670000000e-05,  \
+ 5.645250000000e-05, + 5.669690000000e-05, + 5.693050000000e-05, + 5.715420000000e-05, + 5.736870000000e-05,  \
+ 5.757440000000e-05, + 5.777200000000e-05, + 5.796210000000e-05, + 5.814510000000e-05, + 5.832150000000e-05,  \
+ 5.849170000000e-05, + 5.865610000000e-05, + 5.881510000000e-05, + 5.896900000000e-05, + 5.911820000000e-05,  \
+ 5.926280000000e-05, + 5.940320000000e-05, + 5.953960000000e-05, + 5.967230000000e-05, + 5.980150000000e-05,  \
+ 5.992730000000e-05, + 6.005000000000e-05, + 6.016970000000e-05, + 6.028660000000e-05, + 6.040080000000e-05,  \
+ 6.051240000000e-05, + 6.062170000000e-05, + 6.072870000000e-05, + 6.083360000000e-05, + 6.093630000000e-05 ]

.param id_pred_data_vg0.72=[ \
+ 2.316530444659e-06, + 4.593307676259e-06, + 6.828569748905e-06, + 9.020622237585e-06, + 1.116779603763e-05,  \
+ 1.326848723693e-05, + 1.532113543362e-05, + 1.732428558171e-05, + 1.927648481796e-05, + 2.117643889505e-05,  \
+ 2.302298322320e-05, + 2.481485134922e-05, + 2.655112257344e-05, + 2.823081362294e-05, + 2.985322862514e-05,  \
+ 3.141763852909e-05, + 3.292350156698e-05, + 3.437058854615e-05, + 3.575856258976e-05, + 3.708743606694e-05,  \
+ 3.835737879854e-05, + 3.956862346968e-05, + 4.072166615515e-05, + 4.181723808870e-05, + 4.285612521926e-05,  \
+ 4.383946652524e-05, + 4.476839967538e-05, + 4.564446688164e-05, + 4.646909801522e-05, + 4.724408208858e-05,  \
+ 4.797134955879e-05, + 4.865300375968e-05, + 4.929116723360e-05, + 4.988828004571e-05, + 5.044654317317e-05,  \
+ 5.096858250909e-05, + 5.145687653567e-05, + 5.191398580791e-05, + 5.234257550910e-05, + 5.274498835206e-05,  \
+ 5.312380977557e-05, + 5.348157661501e-05, + 5.382052258938e-05, + 5.414280924015e-05, + 5.445062088256e-05,  \
+ 5.474598277942e-05, + 5.503042237251e-05, + 5.530574591830e-05, + 5.557311145822e-05, + 5.583383972407e-05,  \
+ 5.608892017335e-05, + 5.633913737256e-05, + 5.658507645421e-05, + 5.682708753739e-05, + 5.706552765332e-05,  \
+ 5.730028089602e-05, + 5.753148281656e-05, + 5.775872108643e-05, + 5.798189733468e-05, + 5.820036894875e-05,  \
+ 5.841385216627e-05, + 5.862175763468e-05, + 5.882345256396e-05, + 5.901845637709e-05, + 5.920614348724e-05,  \
+ 5.938597387285e-05, + 5.955744767562e-05, + 5.972021288471e-05, + 5.987361444568e-05, + 6.001737419865e-05,  \
+ 6.015120961820e-05, + 6.027482100762e-05, + 6.038818544766e-05, + 6.049105097190e-05, + 6.058348481019e-05,  \
+ 6.066532747354e-05, + 6.073682321585e-05, + 6.079809187213e-05, + 6.084918444685e-05, + 6.089039379731e-05 ]

* Data table for Id-Vd at Vg = 0.73V
.param vd_data_vg0.73=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.73=[ \
+ 2.306100000000e-06, + 4.593300000000e-06, + 6.854800000000e-06, + 9.084400000000e-06, + 1.127640000000e-05,  \
+ 1.342540000000e-05, + 1.552670000000e-05, + 1.757640000000e-05, + 1.957120000000e-05, + 2.150830000000e-05,  \
+ 2.338550000000e-05, + 2.520120000000e-05, + 2.695420000000e-05, + 2.864380000000e-05, + 3.026940000000e-05,  \
+ 3.183100000000e-05, + 3.332910000000e-05, + 3.476410000000e-05, + 3.613700000000e-05, + 3.744880000000e-05,  \
+ 3.870110000000e-05, + 3.989520000000e-05, + 4.103310000000e-05, + 4.211650000000e-05, + 4.314740000000e-05,  \
+ 4.412790000000e-05, + 4.505990000000e-05, + 4.594540000000e-05, + 4.678660000000e-05, + 4.758520000000e-05,  \
+ 4.834310000000e-05, + 4.906230000000e-05, + 4.974440000000e-05, + 5.039120000000e-05, + 5.100430000000e-05,  \
+ 5.158530000000e-05, + 5.213580000000e-05, + 5.265740000000e-05, + 5.315160000000e-05, + 5.361980000000e-05,  \
+ 5.406350000000e-05, + 5.448410000000e-05, + 5.488300000000e-05, + 5.526130000000e-05, + 5.562050000000e-05,  \
+ 5.596170000000e-05, + 5.628610000000e-05, + 5.659460000000e-05, + 5.688850000000e-05, + 5.716850000000e-05,  \
+ 5.743570000000e-05, + 5.769090000000e-05, + 5.793490000000e-05, + 5.816850000000e-05, + 5.839220000000e-05,  \
+ 5.860690000000e-05, + 5.881300000000e-05, + 5.901110000000e-05, + 5.920180000000e-05, + 5.938550000000e-05,  \
+ 5.956270000000e-05, + 5.973380000000e-05, + 5.989920000000e-05, + 6.005910000000e-05, + 6.021400000000e-05,  \
+ 6.036420000000e-05, + 6.050990000000e-05, + 6.065140000000e-05, + 6.078890000000e-05, + 6.092270000000e-05,  \
+ 6.105290000000e-05, + 6.117980000000e-05, + 6.130360000000e-05, + 6.142440000000e-05, + 6.154240000000e-05,  \
+ 6.165770000000e-05, + 6.177050000000e-05, + 6.188080000000e-05, + 6.198890000000e-05, + 6.209480000000e-05 ]

.param id_pred_data_vg0.73=[ \
+ 2.326384565094e-06, + 4.613730998244e-06, + 6.860331923235e-06, + 9.064507903531e-06, + 1.122467510868e-05,  \
+ 1.333916938165e-05, + 1.540652854601e-05, + 1.742531196214e-05, + 1.939409208717e-05, + 2.131151122740e-05,  \
+ 2.317644175491e-05, + 2.498771063983e-05, + 2.674423609278e-05, + 2.844512404408e-05, + 3.008955027326e-05,  \
+ 3.167682560161e-05, + 3.320641568280e-05, + 3.467790840659e-05, + 3.609102641349e-05, + 3.744560526684e-05,  \
+ 3.874177768012e-05, + 3.997972438810e-05, + 4.115989111597e-05, + 4.228273755871e-05, + 4.334918412496e-05,  \
+ 4.435995477252e-05, + 4.531642291113e-05, + 4.621965286788e-05, + 4.707123662229e-05, + 4.787274228875e-05,  \
+ 4.862600850174e-05, + 4.933309741318e-05, + 4.999591372325e-05, + 5.061676725745e-05, + 5.119787747390e-05,  \
+ 5.174175021239e-05, + 5.225085886195e-05, + 5.272779031657e-05, + 5.317486182321e-05, + 5.359476199374e-05,  \
+ 5.398998313467e-05, + 5.436291714432e-05, + 5.471600816236e-05, + 5.505136621650e-05, + 5.537131728488e-05,  \
+ 5.567772750510e-05, + 5.597256000328e-05, + 5.625742720440e-05, + 5.653370273649e-05, + 5.680284084519e-05,  \
+ 5.706593903597e-05, + 5.732373974752e-05, + 5.757694445492e-05, + 5.782622873085e-05, + 5.807163033751e-05,  \
+ 5.831358139403e-05, + 5.855182957021e-05, + 5.878635100089e-05, + 5.901681775867e-05, + 5.924297729507e-05,  \
+ 5.946408185991e-05, + 5.967987977783e-05, + 5.988972559862e-05, + 6.009296514094e-05, + 6.028912721376e-05,  \
+ 6.047755610780e-05, + 6.065767658583e-05, + 6.082901614718e-05, + 6.099107755290e-05, + 6.114329589764e-05,  \
+ 6.128566332336e-05, + 6.141769874375e-05, + 6.153902242659e-05, + 6.164978112793e-05, + 6.174975897011e-05,  \
+ 6.183890160173e-05, + 6.191727290570e-05, + 6.198499031598e-05, + 6.204222918313e-05, + 6.208915729076e-05 ]

* Data table for Id-Vd at Vg = 0.74V
.param vd_data_vg0.74=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.74=[ \
+ 2.318500000000e-06, + 4.618600000000e-06, + 6.893700000000e-06, + 9.137500000000e-06, + 1.134440000000e-05,  \
+ 1.350900000000e-05, + 1.562680000000e-05, + 1.769370000000e-05, + 1.970640000000e-05, + 2.166220000000e-05,  \
+ 2.355870000000e-05, + 2.539450000000e-05, + 2.716810000000e-05, + 2.887890000000e-05, + 3.052620000000e-05,  \
+ 3.211020000000e-05, + 3.363090000000e-05, + 3.508890000000e-05, + 3.648500000000e-05, + 3.782030000000e-05,  \
+ 3.909600000000e-05, + 4.031380000000e-05, + 4.147510000000e-05, + 4.258190000000e-05, + 4.363600000000e-05,  \
+ 4.463940000000e-05, + 4.559410000000e-05, + 4.650200000000e-05, + 4.736520000000e-05, + 4.818550000000e-05,  \
+ 4.896490000000e-05, + 4.970510000000e-05, + 5.040790000000e-05, + 5.107500000000e-05, + 5.170800000000e-05,  \
+ 5.230860000000e-05, + 5.287820000000e-05, + 5.341850000000e-05, + 5.393090000000e-05, + 5.441680000000e-05,  \
+ 5.487770000000e-05, + 5.531490000000e-05, + 5.572980000000e-05, + 5.612370000000e-05, + 5.649780000000e-05,  \
+ 5.685330000000e-05, + 5.719140000000e-05, + 5.751310000000e-05, + 5.781950000000e-05, + 5.811160000000e-05,  \
+ 5.839030000000e-05, + 5.865640000000e-05, + 5.891090000000e-05, + 5.915440000000e-05, + 5.938760000000e-05,  \
+ 5.961130000000e-05, + 5.982600000000e-05, + 6.003240000000e-05, + 6.023090000000e-05, + 6.042200000000e-05,  \
+ 6.060640000000e-05, + 6.078420000000e-05, + 6.095600000000e-05, + 6.112220000000e-05, + 6.128300000000e-05,  \
+ 6.143880000000e-05, + 6.158980000000e-05, + 6.173650000000e-05, + 6.187900000000e-05, + 6.201750000000e-05,  \
+ 6.215230000000e-05, + 6.228350000000e-05, + 6.241150000000e-05, + 6.253630000000e-05, + 6.265810000000e-05,  \
+ 6.277710000000e-05, + 6.289340000000e-05, + 6.300720000000e-05, + 6.311850000000e-05, + 6.322760000000e-05 ]

.param id_pred_data_vg0.74=[ \
+ 2.335485332878e-06, + 4.632619093172e-06, + 6.889737996971e-06, + 9.105193894356e-06, + 1.127743380493e-05,  \
+ 1.340487040579e-05, + 1.548602987896e-05, + 1.751944073476e-05, + 1.950374833541e-05, + 2.143770980183e-05,  \
+ 2.332002230105e-05, + 2.514956169762e-05, + 2.692529538763e-05, + 2.864633075660e-05, + 3.031175365322e-05,  \
+ 3.192088566720e-05, + 3.347314603161e-05, + 3.496806108160e-05, + 3.640525595983e-05, + 3.778467071243e-05,  \
+ 3.910619096132e-05, + 4.036998405354e-05, + 4.157642120845e-05, + 4.272586433217e-05, + 4.381898907013e-05,  \
+ 4.485675453907e-05, + 4.584006266668e-05, + 4.677004937548e-05, + 4.764822369907e-05, + 4.847586824326e-05,  \
+ 4.925496774376e-05, + 4.998712334782e-05, + 5.067447898909e-05, + 5.131907644682e-05, + 5.192315002205e-05,  \
+ 5.248909641523e-05, + 5.301920697093e-05, + 5.351595900720e-05, + 5.398196706665e-05, + 5.441960529424e-05,  \
+ 5.483146800543e-05, + 5.521990213310e-05, + 5.558735923842e-05, + 5.593621986918e-05, + 5.626844940707e-05,  \
+ 5.658624781063e-05, + 5.689164201613e-05, + 5.718620144762e-05, + 5.747164417699e-05, + 5.774921373813e-05,  \
+ 5.802028899780e-05, + 5.828556924826e-05, + 5.854609524249e-05, + 5.880238124519e-05, + 5.905479483772e-05,  \
+ 5.930361221544e-05, + 5.954886022664e-05, + 5.979034016491e-05, + 6.002800750139e-05, + 6.026148766978e-05,  \
+ 6.049020252249e-05, + 6.071377283661e-05, + 6.093161711760e-05, + 6.114311050624e-05, + 6.134756076790e-05,  \
+ 6.154446018627e-05, + 6.173317517096e-05, + 6.191316031618e-05, + 6.208403603523e-05, + 6.224509124877e-05,  \
+ 6.239603346330e-05, + 6.253648374695e-05, + 6.266623408010e-05, + 6.278519227635e-05, + 6.289294469752e-05,  \
+ 6.298974301899e-05, + 6.307540788839e-05, + 6.315005608485e-05, + 6.321379361907e-05, + 6.326685543172e-05 ]

* Data table for Id-Vd at Vg = 0.75V
.param vd_data_vg0.75=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.75=[ \
+ 2.330500000000e-06, + 4.642900000000e-06, + 6.931000000000e-06, + 9.188500000000e-06, + 1.140980000000e-05,  \
+ 1.358940000000e-05, + 1.572300000000e-05, + 1.780640000000e-05, + 1.983630000000e-05, + 2.180990000000e-05,  \
+ 2.372510000000e-05, + 2.558000000000e-05, + 2.737350000000e-05, + 2.910460000000e-05, + 3.077290000000e-05,  \
+ 3.237810000000e-05, + 3.392060000000e-05, + 3.540060000000e-05, + 3.681910000000e-05, + 3.817690000000e-05,  \
+ 3.947530000000e-05, + 4.071580000000e-05, + 4.189980000000e-05, + 4.302910000000e-05, + 4.410560000000e-05,  \
+ 4.513120000000e-05, + 4.610770000000e-05, + 4.703730000000e-05, + 4.792180000000e-05, + 4.876310000000e-05,  \
+ 4.956320000000e-05, + 5.032380000000e-05, + 5.104660000000e-05, + 5.173340000000e-05, + 5.238590000000e-05,  \
+ 5.300540000000e-05, + 5.359370000000e-05, + 5.415220000000e-05, + 5.468240000000e-05, + 5.518570000000e-05,  \
+ 5.566350000000e-05, + 5.611710000000e-05, + 5.654780000000e-05, + 5.695710000000e-05, + 5.734590000000e-05,  \
+ 5.771570000000e-05, + 5.806750000000e-05, + 5.840230000000e-05, + 5.872130000000e-05, + 5.902550000000e-05,  \
+ 5.931570000000e-05, + 5.959290000000e-05, + 5.985790000000e-05, + 6.011140000000e-05, + 6.035420000000e-05,  \
+ 6.058700000000e-05, + 6.081050000000e-05, + 6.102520000000e-05, + 6.123160000000e-05, + 6.143040000000e-05,  \
+ 6.162190000000e-05, + 6.180670000000e-05, + 6.198500000000e-05, + 6.215750000000e-05, + 6.232430000000e-05,  \
+ 6.248580000000e-05, + 6.264240000000e-05, + 6.279430000000e-05, + 6.294180000000e-05, + 6.308510000000e-05,  \
+ 6.322450000000e-05, + 6.336020000000e-05, + 6.349240000000e-05, + 6.362130000000e-05, + 6.374700000000e-05,  \
+ 6.386980000000e-05, + 6.398970000000e-05, + 6.410690000000e-05, + 6.422160000000e-05, + 6.433390000000e-05 ]

.param id_pred_data_vg0.75=[ \
+ 2.343859378016e-06, + 4.650023474824e-06, + 6.916875281604e-06, + 9.142809431069e-06, + 1.132628094638e-05,  \
+ 1.346574397758e-05, + 1.555976676173e-05, + 1.760693965480e-05, + 1.960590670933e-05, + 2.155532274628e-05,  \
+ 2.345404340304e-05, + 2.530090219807e-05, + 2.709489257541e-05, + 2.883498789743e-05, + 3.052043030038e-05,  \
+ 3.215041942894e-05, + 3.372425911948e-05, + 3.524161234964e-05, + 3.670205303933e-05, + 3.810521448031e-05,  \
+ 3.945114731323e-05, + 4.073995951330e-05, + 4.197177855531e-05, + 4.314704448916e-05, + 4.426626765053e-05,  \
+ 4.533027065918e-05, + 4.633982185624e-05, + 4.729609237984e-05, + 4.820041373023e-05, + 4.905397508992e-05,  \
+ 4.985848441720e-05, + 5.061563104391e-05, + 5.132743928698e-05, + 5.199581122724e-05, + 5.262285485514e-05,  \
+ 5.321073636878e-05, + 5.376202854677e-05, + 5.427893425804e-05, + 5.476401609485e-05, + 5.521962884814e-05,  \
+ 5.564843144384e-05, + 5.605264770566e-05, + 5.643473850796e-05, + 5.679721012712e-05, + 5.714206636185e-05,  \
+ 5.747165414505e-05, + 5.778771970654e-05, + 5.809223977849e-05, + 5.838682525791e-05, + 5.867306390428e-05,  \
+ 5.895207767026e-05, + 5.922494747210e-05, + 5.949273705482e-05, + 5.975590262096e-05, + 6.001521323924e-05,  \
+ 6.027066672686e-05, + 6.052268261556e-05, + 6.077106838347e-05, + 6.101565544668e-05, + 6.125619256636e-05,  \
+ 6.149237837235e-05, + 6.172347741085e-05, + 6.194907669851e-05, + 6.216849200428e-05, + 6.238130699785e-05,  \
+ 6.258665729547e-05, + 6.278395805566e-05, + 6.297265528701e-05, + 6.315228907624e-05, + 6.332215925795e-05,  \
+ 6.348188609991e-05, + 6.363109219819e-05, + 6.376943798386e-05, + 6.389676753315e-05, + 6.401277460100e-05,  \
+ 6.411747570382e-05, + 6.421073514502e-05, + 6.429273300455e-05, + 6.436345815018e-05, + 6.442307494581e-05 ]

* Data table for Id-Vd at Vg = 0.76V
.param vd_data_vg0.76=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.76=[ \
+ 2.341900000000e-06, + 4.666400000000e-06, + 6.967000000000e-06, + 9.237600000000e-06, + 1.147260000000e-05,  \
+ 1.366670000000e-05, + 1.581540000000e-05, + 1.791470000000e-05, + 1.996110000000e-05, + 2.195190000000e-05,  \
+ 2.388490000000e-05, + 2.575830000000e-05, + 2.757070000000e-05, + 2.932140000000e-05, + 3.100960000000e-05,  \
+ 3.263540000000e-05, + 3.419870000000e-05, + 3.569990000000e-05, + 3.713980000000e-05, + 3.851930000000e-05,  \
+ 3.983950000000e-05, + 4.110180000000e-05, + 4.230760000000e-05, + 4.345860000000e-05, + 4.455670000000e-05,  \
+ 4.560370000000e-05, + 4.660140000000e-05, + 4.755190000000e-05, + 4.845700000000e-05, + 4.931860000000e-05,  \
+ 5.013870000000e-05, + 5.091900000000e-05, + 5.166120000000e-05, + 5.236710000000e-05, + 5.303830000000e-05,  \
+ 5.367630000000e-05, + 5.428270000000e-05, + 5.485900000000e-05, + 5.540650000000e-05, + 5.592670000000e-05,  \
+ 5.642100000000e-05, + 5.689070000000e-05, + 5.733710000000e-05, + 5.776140000000e-05, + 5.816490000000e-05,  \
+ 5.854880000000e-05, + 5.891420000000e-05, + 5.926210000000e-05, + 5.959370000000e-05, + 5.990990000000e-05,  \
+ 6.021170000000e-05, + 6.049990000000e-05, + 6.077550000000e-05, + 6.103910000000e-05, + 6.129160000000e-05,  \
+ 6.153370000000e-05, + 6.176590000000e-05, + 6.198900000000e-05, + 6.220350000000e-05, + 6.240990000000e-05,  \
+ 6.260880000000e-05, + 6.280050000000e-05, + 6.298560000000e-05, + 6.316440000000e-05, + 6.333730000000e-05,  \
+ 6.350470000000e-05, + 6.366680000000e-05, + 6.382410000000e-05, + 6.397670000000e-05, + 6.412490000000e-05,  \
+ 6.426900000000e-05, + 6.440920000000e-05, + 6.454570000000e-05, + 6.467880000000e-05, + 6.480850000000e-05,  \
+ 6.493500000000e-05, + 6.505860000000e-05, + 6.517940000000e-05, + 6.529750000000e-05, + 6.541310000000e-05 ]

.param id_pred_data_vg0.76=[ \
+ 2.351536677452e-06, + 4.666011082008e-06, + 6.941835017642e-06, + 9.177447063848e-06, + 1.137135914178e-05,  \
+ 1.352204504656e-05, + 1.562808654853e-05, + 1.768811140209e-05, + 1.970074532437e-05, + 2.166475605918e-05,  \
+ 2.357891804422e-05, + 2.544218266848e-05, + 2.725338898017e-05, + 2.901163126808e-05, + 3.071603860008e-05,  \
+ 3.236585529521e-05, + 3.396044514375e-05, + 3.549922228558e-05, + 3.698183514643e-05, + 3.840795834549e-05,  \
+ 3.977744432632e-05, + 4.109035508009e-05, + 4.234673964675e-05, + 4.354703938588e-05, + 4.469167834031e-05,  \
+ 4.578114254400e-05, + 4.681644699303e-05, + 4.779850714840e-05, + 4.872837220319e-05, + 4.960746009601e-05,  \
+ 5.043710887549e-05, + 5.121911410242e-05, + 5.195511155762e-05, + 5.264706560411e-05, + 5.329695632099e-05,  \
+ 5.390712060034e-05, + 5.447954972624e-05, + 5.501678795554e-05, + 5.552111673751e-05, + 5.599504220299e-05,  \
+ 5.644095101161e-05, + 5.686122720363e-05, + 5.725838374929e-05, + 5.763471475802e-05, + 5.799257414765e-05,  \
+ 5.833395989612e-05, + 5.866102903383e-05, + 5.897572031245e-05, + 5.927959180553e-05, + 5.957452958683e-05,  \
+ 5.986159449094e-05, + 6.014205981046e-05, + 6.041704727977e-05, + 6.068719361792e-05, + 6.095310563978e-05,  \
+ 6.121523794718e-05, + 6.147372390842e-05, + 6.172871711897e-05, + 6.198011789820e-05, + 6.222754163900e-05,  \
+ 6.247074699786e-05, + 6.270923709963e-05, + 6.294240229181e-05, + 6.316972896457e-05, + 6.339056453726e-05,  \
+ 6.360427229083e-05, + 6.381001549016e-05, + 6.400753074558e-05, + 6.419581659429e-05, + 6.437450501835e-05,  \
+ 6.454316440795e-05, + 6.470115738921e-05, + 6.484832607384e-05, + 6.498431306682e-05, + 6.510875755339e-05,  \
+ 6.522171257529e-05, + 6.532299696119e-05, + 6.541265218402e-05, + 6.549067096785e-05, + 6.555726868100e-05 ]

* Data table for Id-Vd at Vg = 0.77V
.param vd_data_vg0.77=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.77=[ \
+ 2.353000000000e-06, + 4.688900000000e-06, + 7.001500000000e-06, + 9.284800000000e-06, + 1.153300000000e-05,  \
+ 1.374110000000e-05, + 1.590430000000e-05, + 1.801870000000e-05, + 2.008100000000e-05, + 2.208840000000e-05,  \
+ 2.403840000000e-05, + 2.592950000000e-05, + 2.776020000000e-05, + 2.952950000000e-05, + 3.123700000000e-05,  \
+ 3.288240000000e-05, + 3.446570000000e-05, + 3.598730000000e-05, + 3.744770000000e-05, + 3.884800000000e-05,  \
+ 4.018910000000e-05, + 4.147230000000e-05, + 4.269910000000e-05, + 4.387110000000e-05, + 4.499000000000e-05,  \
+ 4.605750000000e-05, + 4.707570000000e-05, + 4.804630000000e-05, + 4.897130000000e-05, + 4.985250000000e-05,  \
+ 5.069190000000e-05, + 5.149120000000e-05, + 5.225220000000e-05, + 5.297650000000e-05, + 5.366590000000e-05,  \
+ 5.432170000000e-05, + 5.494560000000e-05, + 5.553910000000e-05, + 5.610350000000e-05, + 5.664020000000e-05,  \
+ 5.715060000000e-05, + 5.763600000000e-05, + 5.809770000000e-05, + 5.853690000000e-05, + 5.895480000000e-05,  \
+ 5.935260000000e-05, + 5.973140000000e-05, + 6.009230000000e-05, + 6.043640000000e-05, + 6.076460000000e-05,  \
+ 6.107790000000e-05, + 6.137720000000e-05, + 6.166330000000e-05, + 6.193710000000e-05, + 6.219930000000e-05,  \
+ 6.245070000000e-05, + 6.269180000000e-05, + 6.292340000000e-05, + 6.314600000000e-05, + 6.336010000000e-05,  \
+ 6.356640000000e-05, + 6.376520000000e-05, + 6.395710000000e-05, + 6.414230000000e-05, + 6.432140000000e-05,  \
+ 6.449470000000e-05, + 6.466250000000e-05, + 6.482520000000e-05, + 6.498300000000e-05, + 6.513620000000e-05,  \
+ 6.528510000000e-05, + 6.542980000000e-05, + 6.557070000000e-05, + 6.570790000000e-05, + 6.584170000000e-05,  \
+ 6.597220000000e-05, + 6.609950000000e-05, + 6.622390000000e-05, + 6.634540000000e-05, + 6.646430000000e-05 ]

.param id_pred_data_vg0.77=[ \
+ 2.358541823924e-06, + 4.680624988396e-06, + 6.964712374611e-06, + 9.209263953380e-06, + 1.141282846220e-05,  \
+ 1.357392029604e-05, + 1.569113897858e-05, + 1.776316668838e-05, + 1.978864398552e-05, + 2.176633570343e-05,  \
+ 2.369507681578e-05, + 2.557371568400e-05, + 2.740123483818e-05, + 2.917663776316e-05, + 3.089910678682e-05,  \
+ 3.256785683334e-05, + 3.418210981181e-05, + 3.574146190658e-05, + 3.724527137820e-05, + 3.869343781844e-05,  \
+ 4.008556177723e-05, + 4.142175341258e-05, + 4.270199395251e-05, + 4.392647766508e-05, + 4.509566861088e-05,  \
+ 4.621009284165e-05, + 4.727051564259e-05, + 4.827770520933e-05, + 4.923280386720e-05, + 5.013691261411e-05,  \
+ 5.099141402752e-05, + 5.179791245610e-05, + 5.255786556518e-05, + 5.327339371433e-05, + 5.394613690441e-05,  \
+ 5.457830673549e-05, + 5.517212048289e-05, + 5.572974128881e-05, + 5.625358113321e-05, + 5.674599087797e-05,  \
+ 5.720922359615e-05, + 5.764589121100e-05, + 5.805838256492e-05, + 5.844894505572e-05, + 5.881993347430e-05,  \
+ 5.917352653341e-05, + 5.951177518000e-05, + 5.983684910461e-05, + 6.015026825480e-05, + 6.045391273801e-05,  \
+ 6.074909921153e-05, + 6.103727326263e-05, + 6.131933827419e-05, + 6.159633674542e-05, + 6.186882819748e-05,  \
+ 6.213738699444e-05, + 6.240232418349e-05, + 6.266374213737e-05, + 6.292164813203e-05, + 6.317578372546e-05,  \
+ 6.342572116409e-05, + 6.367137670168e-05, + 6.391195602191e-05, + 6.414688657969e-05, + 6.437556039600e-05,  \
+ 6.459739161073e-05, + 6.481160096882e-05, + 6.501761352411e-05, + 6.521471397718e-05, + 6.540229151142e-05,  \
+ 6.557977023476e-05, + 6.574682076462e-05, + 6.590290366148e-05, + 6.604759197216e-05, + 6.618088264077e-05,  \
+ 6.630221585510e-05, + 6.641182357271e-05, + 6.650944473222e-05, + 6.659518490778e-05, + 6.666907574981e-05 ]

* Data table for Id-Vd at Vg = 0.78V
.param vd_data_vg0.78=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.78=[ \
+ 2.363600000000e-06, + 4.710600000000e-06, + 7.034800000000e-06, + 9.330200000000e-06, + 1.159120000000e-05,  \
+ 1.381250000000e-05, + 1.598980000000e-05, + 1.811880000000e-05, + 2.019630000000e-05, + 2.221950000000e-05,  \
+ 2.418600000000e-05, + 2.609400000000e-05, + 2.794220000000e-05, + 2.972950000000e-05, + 3.145540000000e-05,  \
+ 3.311950000000e-05, + 3.472200000000e-05, + 3.626310000000e-05, + 3.774330000000e-05, + 3.916350000000e-05,  \
+ 4.052460000000e-05, + 4.182800000000e-05, + 4.307490000000e-05, + 4.426700000000e-05, + 4.540590000000e-05,  \
+ 4.649330000000e-05, + 4.753110000000e-05, + 4.852110000000e-05, + 4.946530000000e-05, + 5.036540000000e-05,  \
+ 5.122340000000e-05, + 5.204110000000e-05, + 5.282010000000e-05, + 5.356220000000e-05, + 5.426900000000e-05,  \
+ 5.494210000000e-05, + 5.558290000000e-05, + 5.619300000000e-05, + 5.677370000000e-05, + 5.732650000000e-05,  \
+ 5.785250000000e-05, + 5.835320000000e-05, + 5.882980000000e-05, + 5.928360000000e-05, + 5.971560000000e-05,  \
+ 6.012710000000e-05, + 6.051920000000e-05, + 6.089290000000e-05, + 6.124940000000e-05, + 6.158950000000e-05,  \
+ 6.191420000000e-05, + 6.222450000000e-05, + 6.252130000000e-05, + 6.280520000000e-05, + 6.307710000000e-05,  \
+ 6.333780000000e-05, + 6.358780000000e-05, + 6.382790000000e-05, + 6.405860000000e-05, + 6.428060000000e-05,  \
+ 6.449430000000e-05, + 6.470030000000e-05, + 6.489890000000e-05, + 6.509070000000e-05, + 6.527610000000e-05,  \
+ 6.545540000000e-05, + 6.562890000000e-05, + 6.579700000000e-05, + 6.596010000000e-05, + 6.611830000000e-05,  \
+ 6.627200000000e-05, + 6.642140000000e-05, + 6.656670000000e-05, + 6.670820000000e-05, + 6.684610000000e-05,  \
+ 6.698050000000e-05, + 6.711160000000e-05, + 6.723960000000e-05, + 6.736470000000e-05, + 6.748690000000e-05 ]

.param id_pred_data_vg0.78=[ \
+ 2.364902320551e-06, + 4.693928058259e-06, + 6.985573272686e-06, + 9.238345082849e-06, + 1.145082278526e-05,  \
+ 1.362157665426e-05, + 1.574921741849e-05, + 1.783241750672e-05, + 1.986990260775e-05, + 2.186044730479e-05,  \
+ 2.380283825914e-05, + 2.569604956079e-05, + 2.753892767942e-05, + 2.933063689852e-05, + 3.107019801973e-05,  \
+ 3.275693161413e-05, + 3.439000269282e-05, + 3.596892056521e-05, + 3.749313313165e-05, + 3.896234265994e-05,  \
+ 4.037626975332e-05, + 4.173488443485e-05, + 4.303806024836e-05, + 4.428602987900e-05, + 4.547914431896e-05,  \
+ 4.661776096327e-05, + 4.770268395077e-05, + 4.873446479905e-05, + 4.971414760803e-05, + 5.064288707217e-05,  \
+ 5.152187804924e-05, + 5.235249176621e-05, + 5.313629197190e-05, + 5.387510231230e-05, + 5.457064107759e-05,  \
+ 5.522497580387e-05, + 5.584015001659e-05, + 5.641823663609e-05, + 5.696164196706e-05, + 5.747263785452e-05,  \
+ 5.795363103971e-05, + 5.840689031174e-05, + 5.883481630008e-05, + 5.923997785430e-05, + 5.962445866317e-05,  \
+ 5.999049462844e-05, + 6.034021120286e-05, + 6.067576585338e-05, + 6.099892591010e-05, + 6.131154077593e-05,  \
+ 6.161496661662e-05, + 6.191073160153e-05, + 6.220009207027e-05, + 6.248381134355e-05, + 6.276292115217e-05,  \
+ 6.303782691248e-05, + 6.330889817036e-05, + 6.357654012390e-05, + 6.384064108715e-05, + 6.410123314708e-05,  \
+ 6.435784234782e-05, + 6.461024808232e-05, + 6.485790290753e-05, + 6.510028615594e-05, + 6.533659252455e-05,  \
+ 6.556642823853e-05, + 6.578886561329e-05, + 6.600326974876e-05, + 6.620898122492e-05, + 6.640543215326e-05,  \
+ 6.659185855824e-05, + 6.676791992504e-05, + 6.693300078041e-05, + 6.708679269650e-05, + 6.722878970322e-05,  \
+ 6.735891365679e-05, + 6.747696286766e-05, + 6.758298011846e-05, + 6.767668382963e-05, + 6.775830406696e-05 ]

* Data table for Id-Vd at Vg = 0.79V
.param vd_data_vg0.79=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.79=[ \
+ 2.373800000000e-06, + 4.731500000000e-06, + 7.066900000000e-06, + 9.373900000000e-06, + 1.164710000000e-05,  \
+ 1.388130000000e-05, + 1.607200000000e-05, + 1.821510000000e-05, + 2.030720000000e-05, + 2.234560000000e-05,  \
+ 2.432780000000e-05, + 2.625210000000e-05, + 2.811700000000e-05, + 2.992160000000e-05, + 3.166510000000e-05,  \
+ 3.334730000000e-05, + 3.496810000000e-05, + 3.652780000000e-05, + 3.802700000000e-05, + 3.946620000000e-05,  \
+ 4.084660000000e-05, + 4.216930000000e-05, + 4.343560000000e-05, + 4.464700000000e-05, + 4.580510000000e-05,  \
+ 4.691150000000e-05, + 4.796820000000e-05, + 4.897690000000e-05, + 4.993950000000e-05, + 5.085790000000e-05,  \
+ 5.173380000000e-05, + 5.256910000000e-05, + 5.336550000000e-05, + 5.412470000000e-05, + 5.484830000000e-05,  \
+ 5.553800000000e-05, + 5.619510000000e-05, + 5.682130000000e-05, + 5.741770000000e-05, + 5.798600000000e-05,  \
+ 5.852720000000e-05, + 5.904280000000e-05, + 5.953390000000e-05, + 6.000180000000e-05, + 6.044760000000e-05,  \
+ 6.087250000000e-05, + 6.127760000000e-05, + 6.166400000000e-05, + 6.203260000000e-05, + 6.238450000000e-05,  \
+ 6.272060000000e-05, + 6.304180000000e-05, + 6.334900000000e-05, + 6.364300000000e-05, + 6.392470000000e-05,  \
+ 6.419460000000e-05, + 6.445350000000e-05, + 6.470220000000e-05, + 6.494110000000e-05, + 6.517090000000e-05,  \
+ 6.539210000000e-05, + 6.560520000000e-05, + 6.581080000000e-05, + 6.600910000000e-05, + 6.620080000000e-05,  \
+ 6.638610000000e-05, + 6.656540000000e-05, + 6.673910000000e-05, + 6.690740000000e-05, + 6.707070000000e-05,  \
+ 6.722930000000e-05, + 6.738340000000e-05, + 6.753320000000e-05, + 6.767900000000e-05, + 6.782100000000e-05,  \
+ 6.795940000000e-05, + 6.809430000000e-05, + 6.822600000000e-05, + 6.835460000000e-05, + 6.848020000000e-05 ]

.param id_pred_data_vg0.79=[ \
+ 2.370651345700e-06, + 4.705985193141e-06, + 7.004532089923e-06, + 9.264849359170e-06, + 1.148552546510e-05,  \
+ 1.366520446027e-05, + 1.580249198014e-05, + 1.789610134438e-05, + 1.994479884161e-05, + 2.194732514909e-05,  \
+ 2.390261055552e-05, + 2.580946544185e-05, + 2.766694233287e-05, + 2.947400556877e-05, + 3.122981215711e-05,  \
+ 3.293356625363e-05, + 3.458457649685e-05, + 3.618215880124e-05, + 3.772591255256e-05, + 3.921538300347e-05,  \
+ 4.065020082635e-05, + 4.203033720842e-05, + 4.335571837146e-05, + 4.462634562515e-05, + 4.584261841956e-05,  \
+ 4.700481280452e-05, + 4.811346661882e-05, + 4.916927486192e-05, + 5.017310395488e-05, + 5.112592043588e-05,  \
+ 5.202902422752e-05, + 5.288349930197e-05, + 5.369086138671e-05, + 5.445280490676e-05, + 5.517100362340e-05,  \
+ 5.584729020484e-05, + 5.648377293255e-05, + 5.708257260267e-05, + 5.764562272816e-05, + 5.817556520924e-05,  \
+ 5.867430460057e-05, + 5.914442619542e-05, + 5.958826688584e-05, + 6.000806286465e-05, + 6.040622174623e-05,  \
+ 6.078505830374e-05, + 6.114646021160e-05, + 6.149288965389e-05, + 6.182594268466e-05, + 6.214765744517e-05,  \
+ 6.245951211895e-05, + 6.276309693931e-05, + 6.305957089353e-05, + 6.335011246847e-05, + 6.363558059093e-05,  \
+ 6.391668401193e-05, + 6.419386059861e-05, + 6.446751620388e-05, + 6.473772780737e-05, + 6.500440067612e-05,  \
+ 6.526742567075e-05, + 6.552633392857e-05, + 6.578088927199e-05, + 6.603030953556e-05, + 6.627410075453e-05,  \
+ 6.651154544670e-05, + 6.674202879367e-05, + 6.696477648802e-05, + 6.717905511323e-05, + 6.738410520484e-05,  \
+ 6.757959985407e-05, + 6.776460155379e-05, + 6.793875552830e-05, + 6.810154911363e-05, + 6.825258788012e-05,  \
+ 6.839167326689e-05, + 6.851845966594e-05, + 6.863298593089e-05, + 6.873496655317e-05, + 6.882474990562e-05 ]

* Data table for Id-Vd at Vg = 0.80V
.param vd_data_vg0.80=[ \
+ 0.010000, + 0.020000, + 0.030000, + 0.040000, + 0.050000, + 0.060000, + 0.070000, + 0.080000, + 0.090000, + 0.100000,  \
+ 0.110000, + 0.120000, + 0.130000, + 0.140000, + 0.150000, + 0.160000, + 0.170000, + 0.180000, + 0.190000, + 0.200000,  \
+ 0.210000, + 0.220000, + 0.230000, + 0.240000, + 0.250000, + 0.260000, + 0.270000, + 0.280000, + 0.290000, + 0.300000,  \
+ 0.310000, + 0.320000, + 0.330000, + 0.340000, + 0.350000, + 0.360000, + 0.370000, + 0.380000, + 0.390000, + 0.400000,  \
+ 0.410000, + 0.420000, + 0.430000, + 0.440000, + 0.450000, + 0.460000, + 0.470000, + 0.480000, + 0.490000, + 0.500000,  \
+ 0.510000, + 0.520000, + 0.530000, + 0.540000, + 0.550000, + 0.560000, + 0.570000, + 0.580000, + 0.590000, + 0.600000,  \
+ 0.610000, + 0.620000, + 0.630000, + 0.640000, + 0.650000, + 0.660000, + 0.670000, + 0.680000, + 0.690000, + 0.700000,  \
+ 0.710000, + 0.720000, + 0.730000, + 0.740000, + 0.750000, + 0.760000, + 0.770000, + 0.780000, + 0.790000, + 0.800000 ]

.param id_actual_data_vg0.80=[ \
+ 2.383700000000e-06, + 4.751600000000e-06, + 7.097700000000e-06, + 9.416100000000e-06, + 1.170100000000e-05,  \
+ 1.394760000000e-05, + 1.615110000000e-05, + 1.830770000000e-05, + 2.041390000000e-05, + 2.246680000000e-05,  \
+ 2.446420000000e-05, + 2.640400000000e-05, + 2.828500000000e-05, + 3.010610000000e-05, + 3.186650000000e-05,  \
+ 3.356600000000e-05, + 3.520440000000e-05, + 3.678200000000e-05, + 3.829920000000e-05, + 3.975680000000e-05,  \
+ 4.115560000000e-05, + 4.249680000000e-05, + 4.378160000000e-05, + 4.501150000000e-05, + 4.618800000000e-05,  \
+ 4.731280000000e-05, + 4.838770000000e-05, + 4.941430000000e-05, + 5.039460000000e-05, + 5.133050000000e-05,  \
+ 5.222360000000e-05, + 5.307580000000e-05, + 5.388890000000e-05, + 5.466460000000e-05, + 5.540440000000e-05,  \
+ 5.611000000000e-05, + 5.678280000000e-05, + 5.742430000000e-05, + 5.803600000000e-05, + 5.861910000000e-05,  \
+ 5.917500000000e-05, + 5.970500000000e-05, + 6.021020000000e-05, + 6.069180000000e-05, + 6.115100000000e-05,  \
+ 6.158900000000e-05, + 6.200680000000e-05, + 6.240550000000e-05, + 6.278610000000e-05, + 6.314960000000e-05,  \
+ 6.349690000000e-05, + 6.382890000000e-05, + 6.414650000000e-05, + 6.445060000000e-05, + 6.474180000000e-05,  \
+ 6.502100000000e-05, + 6.528880000000e-05, + 6.554600000000e-05, + 6.579300000000e-05, + 6.603070000000e-05,  \
+ 6.625940000000e-05, + 6.647970000000e-05, + 6.669210000000e-05, + 6.689710000000e-05, + 6.709510000000e-05,  \
+ 6.728650000000e-05, + 6.747160000000e-05, + 6.765080000000e-05, + 6.782450000000e-05, + 6.799290000000e-05,  \
+ 6.815640000000e-05, + 6.831520000000e-05, + 6.846960000000e-05, + 6.861970000000e-05, + 6.876590000000e-05,  \
+ 6.890830000000e-05, + 6.904710000000e-05, + 6.918250000000e-05, + 6.931460000000e-05, + 6.944370000000e-05 ]

.param id_pred_data_vg0.80=[ \
+ 2.375804906478e-06, + 4.716831608675e-06, + 7.021653873380e-06, + 9.288860601373e-06, + 1.151707037934e-05,  \
+ 1.370497047901e-05, + 1.585118370713e-05, + 1.795449759811e-05, + 2.001362081501e-05, + 2.202742616646e-05,  \
+ 2.399474426056e-05, + 2.591446100269e-05, + 2.778564012260e-05, + 2.960725920275e-05, + 3.137842504657e-05,  \
+ 3.309839870781e-05, + 3.476648926153e-05, + 3.638191003120e-05, + 3.794424555963e-05, + 3.945305943489e-05,  \
+ 4.090799979167e-05, + 4.230891208863e-05, + 4.365565109765e-05, + 4.494822816923e-05, + 4.618688035407e-05,  \
+ 4.737184615806e-05, + 4.850363766309e-05, + 4.958294623066e-05, + 5.061037765699e-05, + 5.158684652997e-05,  \
+ 5.251346156001e-05, + 5.339147057384e-05, + 5.422209724202e-05, + 5.500689730980e-05, + 5.574755050475e-05,  \
+ 5.644592049066e-05, + 5.710366225685e-05, + 5.772306438303e-05, + 5.830600013724e-05, + 5.885475547984e-05,  \
+ 5.937148293015e-05, + 5.985878000502e-05, + 6.031862169039e-05, + 6.075341138057e-05, + 6.116562217358e-05,  \
+ 6.155743845738e-05, + 6.193098728545e-05, + 6.228840211406e-05, + 6.263167510042e-05, + 6.296249921434e-05,  \
+ 6.328296949505e-05, + 6.359438062645e-05, + 6.389825677616e-05, + 6.419553872547e-05, + 6.448752283177e-05,  \
+ 6.477467541117e-05, + 6.505780453153e-05, + 6.533726540511e-05, + 6.561324742506e-05, + 6.588591495529e-05,  \
+ 6.615490165132e-05, + 6.642012143857e-05, + 6.668107096630e-05, + 6.693741772324e-05, + 6.718833574269e-05,  \
+ 6.743317542714e-05, + 6.767149512598e-05, + 6.790226732846e-05, + 6.812487539719e-05, + 6.833874358563e-05,  \
+ 6.854281848064e-05, + 6.873688660562e-05, + 6.892017321661e-05, + 6.909197429195e-05, + 6.925234265509e-05,  \
+ 6.940035091247e-05, + 6.953610107303e-05, + 6.965943946852e-05, + 6.976999284234e-05, + 6.986798834987e-05 ]

* Behavioral voltage sources for Id-Vg plots
EVG_VD0.01 vg_vd0.01 0 VOL='vg_data_vd0.01[min(floor(time*80),79)]'
EID_ACT_VD0.01 id_act_vd0.01 0 VOL='id_actual_data_vd0.01[min(floor(time*80),79)]'
EID_PRED_VD0.01 id_pred_vd0.01 0 VOL='id_pred_data_vd0.01[min(floor(time*80),79)]'

EVG_VD0.20 vg_vd0.20 0 VOL='vg_data_vd0.20[min(floor(time*80),79)]'
EID_ACT_VD0.20 id_act_vd0.20 0 VOL='id_actual_data_vd0.20[min(floor(time*80),79)]'
EID_PRED_VD0.20 id_pred_vd0.20 0 VOL='id_pred_data_vd0.20[min(floor(time*80),79)]'

EVG_VD0.40 vg_vd0.40 0 VOL='vg_data_vd0.40[min(floor(time*80),79)]'
EID_ACT_VD0.40 id_act_vd0.40 0 VOL='id_actual_data_vd0.40[min(floor(time*80),79)]'
EID_PRED_VD0.40 id_pred_vd0.40 0 VOL='id_pred_data_vd0.40[min(floor(time*80),79)]'

EVG_VD0.60 vg_vd0.60 0 VOL='vg_data_vd0.60[min(floor(time*80),79)]'
EID_ACT_VD0.60 id_act_vd0.60 0 VOL='id_actual_data_vd0.60[min(floor(time*80),79)]'
EID_PRED_VD0.60 id_pred_vd0.60 0 VOL='id_pred_data_vd0.60[min(floor(time*80),79)]'

EVG_VD0.80 vg_vd0.80 0 VOL='vg_data_vd0.80[min(floor(time*80),79)]'
EID_ACT_VD0.80 id_act_vd0.80 0 VOL='id_actual_data_vd0.80[min(floor(time*80),79)]'
EID_PRED_VD0.80 id_pred_vd0.80 0 VOL='id_pred_data_vd0.80[min(floor(time*80),79)]'

* Behavioral voltage sources for Id-Vd plots
EVD_VG0.01 vd_vg0.01 0 VOL='vd_data_vg0.01[min(floor(time*80),79)]'
EID_ACT_VG0.01 id_act_vg0.01 0 VOL='id_actual_data_vg0.01[min(floor(time*80),79)]'
EID_PRED_VG0.01 id_pred_vg0.01 0 VOL='id_pred_data_vg0.01[min(floor(time*80),79)]'

EVD_VG0.20 vd_vg0.20 0 VOL='vd_data_vg0.20[min(floor(time*80),79)]'
EID_ACT_VG0.20 id_act_vg0.20 0 VOL='id_actual_data_vg0.20[min(floor(time*80),79)]'
EID_PRED_VG0.20 id_pred_vg0.20 0 VOL='id_pred_data_vg0.20[min(floor(time*80),79)]'

EVD_VG0.40 vd_vg0.40 0 VOL='vd_data_vg0.40[min(floor(time*80),79)]'
EID_ACT_VG0.40 id_act_vg0.40 0 VOL='id_actual_data_vg0.40[min(floor(time*80),79)]'
EID_PRED_VG0.40 id_pred_vg0.40 0 VOL='id_pred_data_vg0.40[min(floor(time*80),79)]'

EVD_VG0.60 vd_vg0.60 0 VOL='vd_data_vg0.60[min(floor(time*80),79)]'
EID_ACT_VG0.60 id_act_vg0.60 0 VOL='id_actual_data_vg0.60[min(floor(time*80),79)]'
EID_PRED_VG0.60 id_pred_vg0.60 0 VOL='id_pred_data_vg0.60[min(floor(time*80),79)]'

EVD_VG0.80 vd_vg0.80 0 VOL='vd_data_vg0.80[min(floor(time*80),79)]'
EID_ACT_VG0.80 id_act_vg0.80 0 VOL='id_actual_data_vg0.80[min(floor(time*80),79)]'
EID_PRED_VG0.80 id_pred_vg0.80 0 VOL='id_pred_data_vg0.80[min(floor(time*80),79)]'

* Run a transient analysis to plot the data
.tran 0.01 1.0

* Plotting hints for WaveView:
* For Id-Vg plots:
*   For Vd=0.01V: Plot V(id_act_vd0.01) vs V(vg_vd0.01) and V(id_pred_vd0.01) vs V(vg_vd0.01)
*   For Vd=0.20V: Plot V(id_act_vd0.20) vs V(vg_vd0.20) and V(id_pred_vd0.20) vs V(vg_vd0.20)
*   For Vd=0.40V: Plot V(id_act_vd0.40) vs V(vg_vd0.40) and V(id_pred_vd0.40) vs V(vg_vd0.40)
*   For Vd=0.60V: Plot V(id_act_vd0.60) vs V(vg_vd0.60) and V(id_pred_vd0.60) vs V(vg_vd0.60)
*   For Vd=0.80V: Plot V(id_act_vd0.80) vs V(vg_vd0.80) and V(id_pred_vd0.80) vs V(vg_vd0.80)
* For Id-Vd plots:
*   For Vg=0.01V: Plot V(id_act_vg0.01) vs V(vd_vg0.01) and V(id_pred_vg0.01) vs V(vd_vg0.01)
*   For Vg=0.20V: Plot V(id_act_vg0.20) vs V(vd_vg0.20) and V(id_pred_vg0.20) vs V(vd_vg0.20)
*   For Vg=0.40V: Plot V(id_act_vg0.40) vs V(vd_vg0.40) and V(id_pred_vg0.40) vs V(vd_vg0.40)
*   For Vg=0.60V: Plot V(id_act_vg0.60) vs V(vd_vg0.60) and V(id_pred_vg0.60) vs V(vd_vg0.60)
*   For Vg=0.80V: Plot V(id_act_vg0.80) vs V(vd_vg0.80) and V(id_pred_vg0.80) vs V(vd_vg0.80)

.end
