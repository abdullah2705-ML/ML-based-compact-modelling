* HSPICE File for IV Comparison - Complete Dataset
* Generated from iv_comparison_sorted.csv

.option abstol=1e-6 reltol=1e-6 post ingold numdgt=8
.hdl "/home/2025_spring/abdullah27/perl5/code/bsimcmg.va"
.include "/home/2025_spring/abdullah27/Research/7nm_FF_160803.pm"

* Parameters
.param vdd = 0.8

******************************************************************
* Original MOSFET Circuit
******************************************************************
* Voltage sources for MOSFET
vd_orig d_orig 0 dc = 0
vg_orig g_orig 0 dc = 0
vs_orig s_orig 0 dc = 0.0
vb_orig b_orig 0 dc = 0

* MOSFET Model (nmos_lvt)
X1 d_orig g_orig s_orig b_orig nmos_lvt L=20n W=100n

******************************************************************
* Common Circuit Components
******************************************************************
* Vd values for our sweep
vd d 0 dc = 0

******************************************************************
* DC Sweeps - One for each selected Vg value
******************************************************************

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.0100) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.0100V
.param vg_value = 0.0100
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.010000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p0100 0 d pwl(0.010000 8.691663e-11 0.020000 1.456779e-10 0.030000 1.861712e-10 
+ 0.040000 2.147540e-10 0.050000 2.355278e-10 0.060000 2.511507e-10 
+ 0.070000 2.633495e-10 0.080000 2.732484e-10 0.090000 2.815800e-10 
+ 0.100000 2.888212e-10 0.110000 2.952821e-10 0.120000 3.011658e-10 
+ 0.130000 3.066067e-10 0.140000 3.116929e-10 0.150000 3.164855e-10 
+ 0.160000 3.210288e-10 0.170000 3.253566e-10 0.180000 3.294980e-10 
+ 0.190000 3.334754e-10 0.200000 3.373139e-10 0.210000 3.410338e-10 
+ 0.220000 3.446564e-10 0.230000 3.482017e-10 0.240000 3.516868e-10 
+ 0.250000 3.551303e-10 0.260000 3.585476e-10 0.270000 3.619549e-10 
+ 0.280000 3.653628e-10 0.290000 3.687843e-10 0.300000 3.722280e-10 
+ 0.310000 3.757040e-10 0.320000 3.792177e-10 0.330000 3.827743e-10 
+ 0.340000 3.863792e-10 0.350000 3.900331e-10 0.360000 3.937402e-10 
+ 0.370000 3.975003e-10 0.380000 4.013137e-10 0.390000 4.051814e-10 
+ 0.400000 4.091013e-10 0.410000 4.130719e-10 0.420000 4.170938e-10 
+ 0.430000 4.211651e-10 0.440000 4.252829e-10 0.450000 4.294451e-10 
+ 0.460000 4.336522e-10 0.470000 4.379007e-10 0.480000 4.421913e-10 
+ 0.490000 4.465209e-10 0.500000 4.508874e-10 0.510000 4.552933e-10 
+ 0.520000 4.597347e-10 0.530000 4.642115e-10 0.540000 4.687251e-10 
+ 0.550000 4.732745e-10 0.560000 4.778606e-10 0.570000 4.824826e-10 
+ 0.580000 4.871414e-10 0.590000 4.918379e-10 0.600000 4.965734e-10 
+ 0.610000 5.013510e-10 0.620000 5.061688e-10 0.630000 5.110306e-10 
+ 0.640000 5.159360e-10 0.650000 5.208905e-10 0.660000 5.258935e-10 
+ 0.670000 5.309481e-10 0.680000 5.360547e-10 0.690000 5.412171e-10 
+ 0.700000 5.464385e-10 0.710000 5.517198e-10 0.720000 5.570627e-10 
+ 0.730000 5.624711e-10 0.740000 5.679468e-10 0.750000 5.734935e-10 
+ 0.760000 5.791108e-10 0.770000 5.848012e-10 0.780000 5.905695e-10 
+ 0.790000 5.964150e-10 0.800000 6.023413e-10)
r_load_0p0100 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.0600) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.0600V
.param vg_value = 0.0600
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.060000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p0600 0 d pwl(0.010000 5.927360e-10 0.020000 9.922707e-10 0.030000 1.263943e-09 
+ 0.040000 1.451069e-09 0.050000 1.582379e-09 0.060000 1.676932e-09 
+ 0.070000 1.747377e-09 0.080000 1.802078e-09 0.090000 1.846567e-09 
+ 0.100000 1.884461e-09 0.110000 1.918110e-09 0.120000 1.949022e-09 
+ 0.130000 1.978142e-09 0.140000 2.006057e-09 0.150000 2.033099e-09 
+ 0.160000 2.059470e-09 0.170000 2.085276e-09 0.180000 2.110559e-09 
+ 0.190000 2.135355e-09 0.200000 2.159691e-09 0.210000 2.183587e-09 
+ 0.220000 2.207069e-09 0.230000 2.230176e-09 0.240000 2.252957e-09 
+ 0.250000 2.275459e-09 0.260000 2.297745e-09 0.270000 2.319886e-09 
+ 0.280000 2.341942e-09 0.290000 2.363978e-09 0.300000 2.386057e-09 
+ 0.310000 2.408243e-09 0.320000 2.430594e-09 0.330000 2.453156e-09 
+ 0.340000 2.475981e-09 0.350000 2.499105e-09 0.360000 2.522555e-09 
+ 0.370000 2.546367e-09 0.380000 2.570561e-09 0.390000 2.595146e-09 
+ 0.400000 2.620133e-09 0.410000 2.645528e-09 0.420000 2.671322e-09 
+ 0.430000 2.697520e-09 0.440000 2.724102e-09 0.450000 2.751046e-09 
+ 0.460000 2.778357e-09 0.470000 2.806005e-09 0.480000 2.833963e-09 
+ 0.490000 2.862203e-09 0.500000 2.890710e-09 0.510000 2.919458e-09 
+ 0.520000 2.948404e-09 0.530000 2.977524e-09 0.540000 3.006796e-09 
+ 0.550000 3.036177e-09 0.560000 3.065644e-09 0.570000 3.095172e-09 
+ 0.580000 3.124714e-09 0.590000 3.154261e-09 0.600000 3.183768e-09 
+ 0.610000 3.213217e-09 0.620000 3.242573e-09 0.630000 3.271814e-09 
+ 0.640000 3.300915e-09 0.650000 3.329856e-09 0.660000 3.358608e-09 
+ 0.670000 3.387153e-09 0.680000 3.415467e-09 0.690000 3.443535e-09 
+ 0.700000 3.471336e-09 0.710000 3.498862e-09 0.720000 3.526094e-09 
+ 0.730000 3.553015e-09 0.740000 3.579620e-09 0.750000 3.605890e-09 
+ 0.760000 3.631831e-09 0.770000 3.657424e-09 0.780000 3.682674e-09 
+ 0.790000 3.707559e-09 0.800000 3.732100e-09)
r_load_0p0600 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.1100) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.1100V
.param vg_value = 0.1100
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.110000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p1100 0 d pwl(0.010000 3.818819e-09 0.020000 6.446108e-09 0.030000 8.259115e-09 
+ 0.040000 9.517726e-09 0.050000 1.040068e-08 0.060000 1.103075e-08 
+ 0.070000 1.149207e-08 0.080000 1.184209e-08 0.090000 1.211990e-08 
+ 0.100000 1.235191e-08 0.110000 1.255568e-08 0.120000 1.274284e-08 
+ 0.130000 1.292070e-08 0.140000 1.309384e-08 0.150000 1.326480e-08 
+ 0.160000 1.343486e-08 0.170000 1.360450e-08 0.180000 1.377352e-08 
+ 0.190000 1.394167e-08 0.200000 1.410836e-08 0.210000 1.427298e-08 
+ 0.220000 1.443506e-08 0.230000 1.459417e-08 0.240000 1.474992e-08 
+ 0.250000 1.490224e-08 0.260000 1.505092e-08 0.270000 1.519607e-08 
+ 0.280000 1.533779e-08 0.290000 1.547641e-08 0.300000 1.561214e-08 
+ 0.310000 1.574538e-08 0.320000 1.587660e-08 0.330000 1.600617e-08 
+ 0.340000 1.613452e-08 0.350000 1.626218e-08 0.360000 1.638946e-08 
+ 0.370000 1.651684e-08 0.380000 1.664473e-08 0.390000 1.677344e-08 
+ 0.400000 1.690331e-08 0.410000 1.703459e-08 0.420000 1.716751e-08 
+ 0.430000 1.730228e-08 0.440000 1.743915e-08 0.450000 1.757808e-08 
+ 0.460000 1.771930e-08 0.470000 1.786282e-08 0.480000 1.800866e-08 
+ 0.490000 1.815681e-08 0.500000 1.830724e-08 0.510000 1.845999e-08 
+ 0.520000 1.861481e-08 0.530000 1.877179e-08 0.540000 1.893071e-08 
+ 0.550000 1.909143e-08 0.560000 1.925397e-08 0.570000 1.941797e-08 
+ 0.580000 1.958338e-08 0.590000 1.975002e-08 0.600000 1.991767e-08 
+ 0.610000 2.008626e-08 0.620000 2.025555e-08 0.630000 2.042528e-08 
+ 0.640000 2.059532e-08 0.650000 2.076551e-08 0.660000 2.093558e-08 
+ 0.670000 2.110551e-08 0.680000 2.127491e-08 0.690000 2.144365e-08 
+ 0.700000 2.161166e-08 0.710000 2.177862e-08 0.720000 2.194445e-08 
+ 0.730000 2.210895e-08 0.740000 2.227196e-08 0.750000 2.243331e-08 
+ 0.760000 2.259284e-08 0.770000 2.275040e-08 0.780000 2.290589e-08 
+ 0.790000 2.305918e-08 0.800000 2.321004e-08)
r_load_0p1100 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.1600) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.1600V
.param vg_value = 0.1600
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.160000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p1600 0 d pwl(0.010000 2.361348e-08 0.020000 4.037383e-08 0.030000 5.224448e-08 
+ 0.040000 6.064482e-08 0.050000 6.659748e-08 0.060000 7.083703e-08 
+ 0.070000 7.388982e-08 0.080000 7.613099e-08 0.090000 7.782761e-08 
+ 0.100000 7.916808e-08 0.110000 8.028476e-08 0.120000 8.126902e-08 
+ 0.130000 8.218355e-08 0.140000 8.306962e-08 0.150000 8.395375e-08 
+ 0.160000 8.485144e-08 0.170000 8.577092e-08 0.180000 8.671494e-08 
+ 0.190000 8.768254e-08 0.200000 8.867026e-08 0.210000 8.967358e-08 
+ 0.220000 9.068683e-08 0.230000 9.170447e-08 0.240000 9.272079e-08 
+ 0.250000 9.373076e-08 0.260000 9.472968e-08 0.270000 9.571384e-08 
+ 0.280000 9.668025e-08 0.290000 9.762659e-08 0.300000 9.855169e-08 
+ 0.310000 9.945465e-08 0.320000 1.003356e-07 0.330000 1.011954e-07 
+ 0.340000 1.020352e-07 0.350000 1.028563e-07 0.360000 1.036614e-07 
+ 0.370000 1.044522e-07 0.380000 1.052311e-07 0.390000 1.060010e-07 
+ 0.400000 1.067639e-07 0.410000 1.075225e-07 0.420000 1.082792e-07 
+ 0.430000 1.090364e-07 0.440000 1.097955e-07 0.450000 1.105594e-07 
+ 0.460000 1.113291e-07 0.470000 1.121063e-07 0.480000 1.128924e-07 
+ 0.490000 1.136885e-07 0.500000 1.144952e-07 0.510000 1.153134e-07 
+ 0.520000 1.161435e-07 0.530000 1.169860e-07 0.540000 1.178408e-07 
+ 0.550000 1.187081e-07 0.560000 1.195874e-07 0.570000 1.204787e-07 
+ 0.580000 1.213817e-07 0.590000 1.222957e-07 0.600000 1.232200e-07 
+ 0.610000 1.241539e-07 0.620000 1.250965e-07 0.630000 1.260474e-07 
+ 0.640000 1.270053e-07 0.650000 1.279694e-07 0.660000 1.289386e-07 
+ 0.670000 1.299117e-07 0.680000 1.308878e-07 0.690000 1.318657e-07 
+ 0.700000 1.328444e-07 0.710000 1.338227e-07 0.720000 1.347995e-07 
+ 0.730000 1.357735e-07 0.740000 1.367433e-07 0.750000 1.377082e-07 
+ 0.760000 1.386667e-07 0.770000 1.396178e-07 0.780000 1.405601e-07 
+ 0.790000 1.414931e-07 0.800000 1.424147e-07)
r_load_0p1600 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.2200) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.2200V
.param vg_value = 0.2200
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.220000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p2200 0 d pwl(0.010000 1.638347e-07 0.020000 2.884578e-07 0.030000 3.828817e-07 
+ 0.040000 4.541664e-07 0.050000 5.078164e-07 0.060000 5.481073e-07 
+ 0.070000 5.783460e-07 0.080000 6.010841e-07 0.090000 6.182780e-07 
+ 0.100000 6.314235e-07 0.110000 6.416612e-07 0.120000 6.498524e-07 
+ 0.130000 6.566435e-07 0.140000 6.625191e-07 0.150000 6.678313e-07 
+ 0.160000 6.728385e-07 0.170000 6.777204e-07 0.180000 6.826001e-07 
+ 0.190000 6.875587e-07 0.200000 6.926427e-07 0.210000 6.978736e-07 
+ 0.220000 7.032543e-07 0.230000 7.087762e-07 0.240000 7.144216e-07 
+ 0.250000 7.201677e-07 0.260000 7.259856e-07 0.270000 7.318496e-07 
+ 0.280000 7.377318e-07 0.290000 7.436058e-07 0.300000 7.494490e-07 
+ 0.310000 7.552417e-07 0.320000 7.609677e-07 0.330000 7.666131e-07 
+ 0.340000 7.721720e-07 0.350000 7.776360e-07 0.360000 7.830047e-07 
+ 0.370000 7.882799e-07 0.380000 7.934644e-07 0.390000 7.985644e-07 
+ 0.400000 8.035888e-07 0.410000 8.085486e-07 0.420000 8.134538e-07 
+ 0.430000 8.183133e-07 0.440000 8.231420e-07 0.450000 8.279512e-07 
+ 0.460000 8.327513e-07 0.470000 8.375539e-07 0.480000 8.423699e-07 
+ 0.490000 8.472069e-07 0.500000 8.520743e-07 0.510000 8.569782e-07 
+ 0.520000 8.619258e-07 0.530000 8.669186e-07 0.540000 8.719633e-07 
+ 0.550000 8.770595e-07 0.560000 8.822083e-07 0.570000 8.874108e-07 
+ 0.580000 8.926645e-07 0.590000 8.979684e-07 0.600000 9.033164e-07 
+ 0.610000 9.087074e-07 0.620000 9.141332e-07 0.630000 9.195907e-07 
+ 0.640000 9.250727e-07 0.650000 9.305714e-07 0.660000 9.360785e-07 
+ 0.670000 9.415896e-07 0.680000 9.470938e-07 0.690000 9.525821e-07 
+ 0.700000 9.580491e-07 0.710000 9.634785e-07 0.720000 9.688703e-07 
+ 0.730000 9.742066e-07 0.740000 9.794855e-07 0.750000 9.846901e-07 
+ 0.760000 9.898182e-07 0.770000 9.948558e-07 0.780000 9.997942e-07 
+ 0.790000 1.004627e-06 0.800000 1.009341e-06)
r_load_0p2200 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.2700) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.2700V
.param vg_value = 0.2700
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.270000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p2700 0 d pwl(0.010000 4.852416e-07 0.020000 8.815071e-07 0.030000 1.204169e-06 
+ 0.040000 1.466181e-06 0.050000 1.678416e-06 0.060000 1.849984e-06 
+ 0.070000 1.988452e-06 0.080000 2.100105e-06 0.090000 2.190153e-06 
+ 0.100000 2.262871e-06 0.110000 2.321784e-06 0.120000 2.369764e-06 
+ 0.130000 2.409151e-06 0.140000 2.441851e-06 0.150000 2.469390e-06 
+ 0.160000 2.493001e-06 0.170000 2.513655e-06 0.180000 2.532133e-06 
+ 0.190000 2.549044e-06 0.200000 2.564863e-06 0.210000 2.579935e-06 
+ 0.220000 2.594537e-06 0.230000 2.608868e-06 0.240000 2.623064e-06 
+ 0.250000 2.637225e-06 0.260000 2.651405e-06 0.270000 2.665640e-06 
+ 0.280000 2.679943e-06 0.290000 2.694307e-06 0.300000 2.708727e-06 
+ 0.310000 2.723176e-06 0.320000 2.737641e-06 0.330000 2.752097e-06 
+ 0.340000 2.766518e-06 0.350000 2.780894e-06 0.360000 2.795202e-06 
+ 0.370000 2.809433e-06 0.380000 2.823579e-06 0.390000 2.837641e-06 
+ 0.400000 2.851611e-06 0.410000 2.865496e-06 0.420000 2.879305e-06 
+ 0.430000 2.893047e-06 0.440000 2.906732e-06 0.450000 2.920373e-06 
+ 0.460000 2.933986e-06 0.470000 2.947588e-06 0.480000 2.961186e-06 
+ 0.490000 2.974794e-06 0.500000 2.988426e-06 0.510000 3.002090e-06 
+ 0.520000 3.015793e-06 0.530000 3.029534e-06 0.540000 3.043329e-06 
+ 0.550000 3.057166e-06 0.560000 3.071051e-06 0.570000 3.084963e-06 
+ 0.580000 3.098906e-06 0.590000 3.112871e-06 0.600000 3.126827e-06 
+ 0.610000 3.140779e-06 0.620000 3.154694e-06 0.630000 3.168553e-06 
+ 0.640000 3.182339e-06 0.650000 3.196023e-06 0.660000 3.209585e-06 
+ 0.670000 3.222997e-06 0.680000 3.236225e-06 0.690000 3.249247e-06 
+ 0.700000 3.262031e-06 0.710000 3.274548e-06 0.720000 3.286774e-06 
+ 0.730000 3.298673e-06 0.740000 3.310215e-06 0.750000 3.321368e-06 
+ 0.760000 3.332113e-06 0.770000 3.342422e-06 0.780000 3.352254e-06 
+ 0.790000 3.361596e-06 0.800000 3.370410e-06)
r_load_0p2700 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.3200) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.3200V
.param vg_value = 0.3200
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.320000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p3200 0 d pwl(0.010000 9.000973e-07 0.020000 1.681072e-06 0.030000 2.356989e-06 
+ 0.040000 2.940545e-06 0.050000 3.443158e-06 0.060000 3.875066e-06 
+ 0.070000 4.245406e-06 0.080000 4.562346e-06 0.090000 4.833095e-06 
+ 0.100000 5.064052e-06 0.110000 5.260852e-06 0.120000 5.428439e-06 
+ 0.130000 5.571147e-06 0.140000 5.692753e-06 0.150000 5.796542e-06 
+ 0.160000 5.885363e-06 0.170000 5.961656e-06 0.180000 6.027548e-06 
+ 0.190000 6.084828e-06 0.200000 6.135043e-06 0.210000 6.179496e-06 
+ 0.220000 6.219301e-06 0.230000 6.255366e-06 0.240000 6.288479e-06 
+ 0.250000 6.319277e-06 0.260000 6.348289e-06 0.270000 6.375947e-06 
+ 0.280000 6.402601e-06 0.290000 6.428530e-06 0.300000 6.453957e-06 
+ 0.310000 6.479054e-06 0.320000 6.503959e-06 0.330000 6.528770e-06 
+ 0.340000 6.553555e-06 0.350000 6.578374e-06 0.360000 6.603248e-06 
+ 0.370000 6.628219e-06 0.380000 6.653283e-06 0.390000 6.678460e-06 
+ 0.400000 6.703733e-06 0.410000 6.729111e-06 0.420000 6.754605e-06 
+ 0.430000 6.780191e-06 0.440000 6.805873e-06 0.450000 6.831634e-06 
+ 0.460000 6.857493e-06 0.470000 6.883426e-06 0.480000 6.909439e-06 
+ 0.490000 6.935528e-06 0.500000 6.961671e-06 0.510000 6.987875e-06 
+ 0.520000 7.014123e-06 0.530000 7.040404e-06 0.540000 7.066713e-06 
+ 0.550000 7.093029e-06 0.560000 7.119315e-06 0.570000 7.145560e-06 
+ 0.580000 7.171738e-06 0.590000 7.197815e-06 0.600000 7.223744e-06 
+ 0.610000 7.249509e-06 0.620000 7.275040e-06 0.630000 7.300308e-06 
+ 0.640000 7.325270e-06 0.650000 7.349869e-06 0.660000 7.374057e-06 
+ 0.670000 7.397761e-06 0.680000 7.420929e-06 0.690000 7.443511e-06 
+ 0.700000 7.465454e-06 0.710000 7.486685e-06 0.720000 7.507144e-06 
+ 0.730000 7.526775e-06 0.740000 7.545515e-06 0.750000 7.563289e-06 
+ 0.760000 7.580060e-06 0.770000 7.595757e-06 0.780000 7.610347e-06 
+ 0.790000 7.623741e-06 0.800000 7.635906e-06)
r_load_0p3200 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.3700) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.3700V
.param vg_value = 0.3700
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.370000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p3700 0 d pwl(0.010000 1.262592e-06 0.020000 2.407824e-06 0.030000 3.443980e-06 
+ 0.040000 4.379052e-06 0.050000 5.220705e-06 0.060000 5.976271e-06 
+ 0.070000 6.652783e-06 0.080000 7.256902e-06 0.090000 7.794951e-06 
+ 0.100000 8.272930e-06 0.110000 8.696480e-06 0.120000 9.070868e-06 
+ 0.130000 9.401065e-06 0.140000 9.691682e-06 0.150000 9.946963e-06 
+ 0.160000 1.017088e-05 0.170000 1.036706e-05 0.180000 1.053885e-05 
+ 0.190000 1.068925e-05 0.200000 1.082103e-05 0.210000 1.093669e-05 
+ 0.220000 1.103846e-05 0.230000 1.112836e-05 0.240000 1.120816e-05 
+ 0.250000 1.127947e-05 0.260000 1.134365e-05 0.270000 1.140194e-05 
+ 0.280000 1.145543e-05 0.290000 1.150501e-05 0.300000 1.155143e-05 
+ 0.310000 1.159542e-05 0.320000 1.163752e-05 0.330000 1.167822e-05 
+ 0.340000 1.171787e-05 0.350000 1.175682e-05 0.360000 1.179531e-05 
+ 0.370000 1.183351e-05 0.380000 1.187162e-05 0.390000 1.190975e-05 
+ 0.400000 1.194796e-05 0.410000 1.198633e-05 0.420000 1.202485e-05 
+ 0.430000 1.206359e-05 0.440000 1.210250e-05 0.450000 1.214161e-05 
+ 0.460000 1.218091e-05 0.470000 1.222034e-05 0.480000 1.225991e-05 
+ 0.490000 1.229959e-05 0.500000 1.233931e-05 0.510000 1.237908e-05 
+ 0.520000 1.241887e-05 0.530000 1.245861e-05 0.540000 1.249826e-05 
+ 0.550000 1.253781e-05 0.560000 1.257721e-05 0.570000 1.261641e-05 
+ 0.580000 1.265534e-05 0.590000 1.269398e-05 0.600000 1.273228e-05 
+ 0.610000 1.277016e-05 0.620000 1.280759e-05 0.630000 1.284449e-05 
+ 0.640000 1.288079e-05 0.650000 1.291643e-05 0.660000 1.295132e-05 
+ 0.670000 1.298541e-05 0.680000 1.301861e-05 0.690000 1.305083e-05 
+ 0.700000 1.308199e-05 0.710000 1.311203e-05 0.720000 1.314084e-05 
+ 0.730000 1.316836e-05 0.740000 1.319447e-05 0.750000 1.321911e-05 
+ 0.760000 1.324218e-05 0.770000 1.326361e-05 0.780000 1.328328e-05 
+ 0.790000 1.330113e-05 0.800000 1.331709e-05)
r_load_0p3700 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.4300) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.4300V
.param vg_value = 0.4300
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.430000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p4300 0 d pwl(0.010000 1.587107e-06 0.020000 3.077285e-06 0.030000 4.472976e-06 
+ 0.040000 5.776833e-06 0.050000 6.991661e-06 0.060000 8.120492e-06 
+ 0.070000 9.166458e-06 0.080000 1.013291e-05 0.090000 1.102326e-05 
+ 0.100000 1.184114e-05 0.110000 1.259019e-05 0.120000 1.327413e-05 
+ 0.130000 1.389675e-05 0.140000 1.446190e-05 0.150000 1.497341e-05 
+ 0.160000 1.543503e-05 0.170000 1.585055e-05 0.180000 1.622360e-05 
+ 0.190000 1.655781e-05 0.200000 1.685663e-05 0.210000 1.712339e-05 
+ 0.220000 1.736126e-05 0.230000 1.757326e-05 0.240000 1.776233e-05 
+ 0.250000 1.793104e-05 0.260000 1.808190e-05 0.270000 1.821725e-05 
+ 0.280000 1.833911e-05 0.290000 1.844945e-05 0.300000 1.855002e-05 
+ 0.310000 1.864236e-05 0.320000 1.872773e-05 0.330000 1.880751e-05 
+ 0.340000 1.888262e-05 0.350000 1.895404e-05 0.360000 1.902250e-05 
+ 0.370000 1.908866e-05 0.380000 1.915303e-05 0.390000 1.921608e-05 
+ 0.400000 1.927813e-05 0.410000 1.933945e-05 0.420000 1.940025e-05 
+ 0.430000 1.946067e-05 0.440000 1.952078e-05 0.450000 1.958064e-05 
+ 0.460000 1.964029e-05 0.470000 1.969968e-05 0.480000 1.975886e-05 
+ 0.490000 1.981770e-05 0.500000 1.987622e-05 0.510000 1.993432e-05 
+ 0.520000 1.999196e-05 0.530000 2.004904e-05 0.540000 2.010554e-05 
+ 0.550000 2.016137e-05 0.560000 2.021647e-05 0.570000 2.027076e-05 
+ 0.580000 2.032426e-05 0.590000 2.037679e-05 0.600000 2.042836e-05 
+ 0.610000 2.047894e-05 0.620000 2.052842e-05 0.630000 2.057677e-05 
+ 0.640000 2.062393e-05 0.650000 2.066985e-05 0.660000 2.071443e-05 
+ 0.670000 2.075763e-05 0.680000 2.079942e-05 0.690000 2.083970e-05 
+ 0.700000 2.087843e-05 0.710000 2.091547e-05 0.720000 2.095083e-05 
+ 0.730000 2.098439e-05 0.740000 2.101607e-05 0.750000 2.104583e-05 
+ 0.760000 2.107354e-05 0.770000 2.109918e-05 0.780000 2.112256e-05 
+ 0.790000 2.114372e-05 0.800000 2.116246e-05)
r_load_0p4300 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.4800) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.4800V
.param vg_value = 0.4800
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.480000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p4800 0 d pwl(0.010000 1.790846e-06 0.020000 3.502264e-06 0.030000 5.134037e-06 
+ 0.040000 6.686165e-06 0.050000 8.158932e-06 0.060000 9.552805e-06 
+ 0.070000 1.086859e-05 0.080000 1.210729e-05 0.090000 1.327022e-05 
+ 0.100000 1.435891e-05 0.110000 1.537516e-05 0.120000 1.632104e-05 
+ 0.130000 1.719879e-05 0.140000 1.801090e-05 0.150000 1.876003e-05 
+ 0.160000 1.944901e-05 0.170000 2.008087e-05 0.180000 2.065864e-05 
+ 0.190000 2.118558e-05 0.200000 2.166485e-05 0.210000 2.209982e-05 
+ 0.220000 2.249372e-05 0.230000 2.284984e-05 0.240000 2.317139e-05 
+ 0.250000 2.346146e-05 0.260000 2.372312e-05 0.270000 2.395930e-05 
+ 0.280000 2.417273e-05 0.290000 2.436601e-05 0.300000 2.454165e-05 
+ 0.310000 2.470194e-05 0.320000 2.484886e-05 0.330000 2.498441e-05 
+ 0.340000 2.511025e-05 0.350000 2.522800e-05 0.360000 2.533892e-05 
+ 0.370000 2.544425e-05 0.380000 2.554498e-05 0.390000 2.564198e-05 
+ 0.400000 2.573598e-05 0.410000 2.582751e-05 0.420000 2.591709e-05 
+ 0.430000 2.600506e-05 0.440000 2.609167e-05 0.450000 2.617712e-05 
+ 0.460000 2.626150e-05 0.470000 2.634485e-05 0.480000 2.642727e-05 
+ 0.490000 2.650859e-05 0.500000 2.658885e-05 0.510000 2.666797e-05 
+ 0.520000 2.674582e-05 0.530000 2.682233e-05 0.540000 2.689739e-05 
+ 0.550000 2.697084e-05 0.560000 2.704264e-05 0.570000 2.711273e-05 
+ 0.580000 2.718097e-05 0.590000 2.724724e-05 0.600000 2.731160e-05 
+ 0.610000 2.737382e-05 0.620000 2.743402e-05 0.630000 2.749202e-05 
+ 0.640000 2.754785e-05 0.650000 2.760145e-05 0.660000 2.765275e-05 
+ 0.670000 2.770183e-05 0.680000 2.774855e-05 0.690000 2.779296e-05 
+ 0.700000 2.783502e-05 0.710000 2.787464e-05 0.720000 2.791190e-05 
+ 0.730000 2.794673e-05 0.740000 2.797911e-05 0.750000 2.800894e-05 
+ 0.760000 2.803626e-05 0.770000 2.806106e-05 0.780000 2.808324e-05 
+ 0.790000 2.810274e-05 0.800000 2.811962e-05)
r_load_0p4800 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.5300) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.5300V
.param vg_value = 0.5300
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.530000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p5300 0 d pwl(0.010000 1.954049e-06 0.020000 3.842467e-06 0.030000 5.663767e-06 
+ 0.040000 7.416645e-06 0.050000 9.100011e-06 0.060000 1.071298e-05 
+ 0.070000 1.225490e-05 0.080000 1.372537e-05 0.090000 1.512420e-05 
+ 0.100000 1.645154e-05 0.110000 1.770774e-05 0.120000 1.889345e-05 
+ 0.130000 2.000964e-05 0.140000 2.105737e-05 0.150000 2.203821e-05 
+ 0.160000 2.295378e-05 0.170000 2.380606e-05 0.180000 2.459719e-05 
+ 0.190000 2.532957e-05 0.200000 2.600573e-05 0.210000 2.662844e-05 
+ 0.220000 2.720046e-05 0.230000 2.772483e-05 0.240000 2.820452e-05 
+ 0.250000 2.864266e-05 0.260000 2.904229e-05 0.270000 2.940655e-05 
+ 0.280000 2.973855e-05 0.290000 3.004118e-05 0.300000 3.031735e-05 
+ 0.310000 3.056990e-05 0.320000 3.080143e-05 0.330000 3.101447e-05 
+ 0.340000 3.121125e-05 0.350000 3.139403e-05 0.360000 3.156473e-05 
+ 0.370000 3.172510e-05 0.380000 3.187676e-05 0.390000 3.202113e-05 
+ 0.400000 3.215939e-05 0.410000 3.229255e-05 0.420000 3.242148e-05 
+ 0.430000 3.254691e-05 0.440000 3.266934e-05 0.450000 3.278928e-05 
+ 0.460000 3.290699e-05 0.470000 3.302268e-05 0.480000 3.313638e-05 
+ 0.490000 3.324821e-05 0.500000 3.335807e-05 0.510000 3.346601e-05 
+ 0.520000 3.357180e-05 0.530000 3.367532e-05 0.540000 3.377645e-05 
+ 0.550000 3.387492e-05 0.560000 3.397073e-05 0.570000 3.406362e-05 
+ 0.580000 3.415339e-05 0.590000 3.423997e-05 0.600000 3.432326e-05 
+ 0.610000 3.440309e-05 0.620000 3.447938e-05 0.630000 3.455201e-05 
+ 0.640000 3.462099e-05 0.650000 3.468631e-05 0.660000 3.474792e-05 
+ 0.670000 3.480581e-05 0.680000 3.485988e-05 0.690000 3.491031e-05 
+ 0.700000 3.495708e-05 0.710000 3.500013e-05 0.720000 3.503963e-05 
+ 0.730000 3.507545e-05 0.740000 3.510780e-05 0.750000 3.513661e-05 
+ 0.760000 3.516200e-05 0.770000 3.518398e-05 0.780000 3.520257e-05 
+ 0.790000 3.521778e-05 0.800000 3.522973e-05)
r_load_0p5300 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.5800) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.5800V
.param vg_value = 0.5800
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.580000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p5800 0 d pwl(0.010000 2.085660e-06 0.020000 4.115762e-06 0.030000 6.088336e-06 
+ 0.040000 8.001575e-06 0.050000 9.853797e-06 0.060000 1.164348e-05 
+ 0.070000 1.336926e-05 0.080000 1.503001e-05 0.090000 1.662468e-05 
+ 0.100000 1.815265e-05 0.110000 1.961328e-05 0.120000 2.100637e-05 
+ 0.130000 2.233180e-05 0.140000 2.358984e-05 0.150000 2.478087e-05 
+ 0.160000 2.590570e-05 0.170000 2.696526e-05 0.180000 2.796074e-05 
+ 0.190000 2.889364e-05 0.200000 2.976565e-05 0.210000 3.057869e-05 
+ 0.220000 3.133499e-05 0.230000 3.203671e-05 0.240000 3.268647e-05 
+ 0.250000 3.328687e-05 0.260000 3.384067e-05 0.270000 3.435080e-05 
+ 0.280000 3.482005e-05 0.290000 3.525140e-05 0.300000 3.564793e-05 
+ 0.310000 3.601251e-05 0.320000 3.634800e-05 0.330000 3.665727e-05 
+ 0.340000 3.694316e-05 0.350000 3.720805e-05 0.360000 3.745453e-05 
+ 0.370000 3.768491e-05 0.380000 3.790123e-05 0.390000 3.810546e-05 
+ 0.400000 3.829942e-05 0.410000 3.848472e-05 0.420000 3.866255e-05 
+ 0.430000 3.883415e-05 0.440000 3.900054e-05 0.450000 3.916243e-05 
+ 0.460000 3.932060e-05 0.470000 3.947536e-05 0.480000 3.962710e-05 
+ 0.490000 3.977612e-05 0.500000 3.992244e-05 0.510000 4.006603e-05 
+ 0.520000 4.020686e-05 0.530000 4.034481e-05 0.540000 4.047963e-05 
+ 0.550000 4.061119e-05 0.560000 4.073911e-05 0.570000 4.086314e-05 
+ 0.580000 4.098313e-05 0.590000 4.109878e-05 0.600000 4.120987e-05 
+ 0.610000 4.131609e-05 0.620000 4.141741e-05 0.630000 4.151357e-05 
+ 0.640000 4.160438e-05 0.650000 4.168983e-05 0.660000 4.176987e-05 
+ 0.670000 4.184431e-05 0.680000 4.191328e-05 0.690000 4.197676e-05 
+ 0.700000 4.203472e-05 0.710000 4.208729e-05 0.720000 4.213446e-05 
+ 0.730000 4.217637e-05 0.740000 4.221309e-05 0.750000 4.224487e-05 
+ 0.760000 4.227157e-05 0.770000 4.229343e-05 0.780000 4.231062e-05 
+ 0.790000 4.232321e-05 0.800000 4.233136e-05)
r_load_0p5800 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.6400) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.6400V
.param vg_value = 0.6400
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.640000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p6400 0 d pwl(0.010000 2.207525e-06 0.020000 4.367905e-06 0.030000 6.479159e-06 
+ 0.040000 8.539340e-06 0.050000 1.054661e-05 0.060000 1.249925e-05 
+ 0.070000 1.439561e-05 0.080000 1.623423e-05 0.090000 1.801371e-05 
+ 0.100000 1.973283e-05 0.110000 2.139055e-05 0.120000 2.298600e-05 
+ 0.130000 2.451843e-05 0.140000 2.598734e-05 0.150000 2.739235e-05 
+ 0.160000 2.873347e-05 0.170000 3.001080e-05 0.180000 3.122457e-05 
+ 0.190000 3.237540e-05 0.200000 3.346406e-05 0.210000 3.449158e-05 
+ 0.220000 3.545914e-05 0.230000 3.636826e-05 0.240000 3.722056e-05 
+ 0.250000 3.801792e-05 0.260000 3.876242e-05 0.270000 3.945620e-05 
+ 0.280000 4.010172e-05 0.290000 4.070138e-05 0.300000 4.125787e-05 
+ 0.310000 4.177390e-05 0.320000 4.225224e-05 0.330000 4.269564e-05 
+ 0.340000 4.310695e-05 0.350000 4.348888e-05 0.360000 4.384424e-05 
+ 0.370000 4.417564e-05 0.380000 4.448568e-05 0.390000 4.477674e-05 
+ 0.400000 4.505116e-05 0.410000 4.531107e-05 0.420000 4.555844e-05 
+ 0.430000 4.579505e-05 0.440000 4.602241e-05 0.450000 4.624211e-05 
+ 0.460000 4.645509e-05 0.470000 4.666253e-05 0.480000 4.686510e-05 
+ 0.490000 4.706346e-05 0.500000 4.725808e-05 0.510000 4.744926e-05 
+ 0.520000 4.763703e-05 0.530000 4.782158e-05 0.540000 4.800267e-05 
+ 0.550000 4.818018e-05 0.560000 4.835380e-05 0.570000 4.852331e-05 
+ 0.580000 4.868831e-05 0.590000 4.884829e-05 0.600000 4.900299e-05 
+ 0.610000 4.915207e-05 0.620000 4.929508e-05 0.630000 4.943153e-05 
+ 0.640000 4.956136e-05 0.650000 4.968418e-05 0.660000 4.979984e-05 
+ 0.670000 4.990797e-05 0.680000 5.000844e-05 0.690000 5.010133e-05 
+ 0.700000 5.018639e-05 0.710000 5.026373e-05 0.720000 5.033327e-05 
+ 0.730000 5.039519e-05 0.740000 5.044946e-05 0.750000 5.049630e-05 
+ 0.760000 5.053588e-05 0.770000 5.056828e-05 0.780000 5.059367e-05 
+ 0.790000 5.061228e-05 0.800000 5.062444e-05)
r_load_0p6400 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.6900) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.6900V
.param vg_value = 0.6900
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.690000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p6900 0 d pwl(0.010000 2.282193e-06 0.020000 4.522242e-06 0.030000 6.718261e-06 
+ 0.040000 8.868465e-06 0.050000 1.097109e-05 0.060000 1.302444e-05 
+ 0.070000 1.502691e-05 0.080000 1.697701e-05 0.090000 1.887326e-05 
+ 0.100000 2.071433e-05 0.110000 2.249903e-05 0.120000 2.422629e-05 
+ 0.130000 2.589509e-05 0.140000 2.750467e-05 0.150000 2.905433e-05 
+ 0.160000 3.054356e-05 0.170000 3.197206e-05 0.180000 3.333956e-05 
+ 0.190000 3.464619e-05 0.200000 3.589218e-05 0.210000 3.707786e-05 
+ 0.220000 3.820375e-05 0.230000 3.927085e-05 0.240000 4.028007e-05 
+ 0.250000 4.123265e-05 0.260000 4.212994e-05 0.270000 4.297352e-05 
+ 0.280000 4.376527e-05 0.290000 4.450703e-05 0.300000 4.520098e-05 
+ 0.310000 4.584916e-05 0.320000 4.645425e-05 0.330000 4.701849e-05 
+ 0.340000 4.754452e-05 0.350000 4.803494e-05 0.360000 4.849242e-05 
+ 0.370000 4.891952e-05 0.380000 4.931903e-05 0.390000 4.969344e-05 
+ 0.400000 5.004536e-05 0.410000 5.037711e-05 0.420000 5.069105e-05 
+ 0.430000 5.098940e-05 0.440000 5.127419e-05 0.450000 5.154740e-05 
+ 0.460000 5.181041e-05 0.470000 5.206495e-05 0.480000 5.231222e-05 
+ 0.490000 5.255328e-05 0.500000 5.278917e-05 0.510000 5.302048e-05 
+ 0.520000 5.324766e-05 0.530000 5.347103e-05 0.540000 5.369091e-05 
+ 0.550000 5.390730e-05 0.560000 5.411997e-05 0.570000 5.432870e-05 
+ 0.580000 5.453331e-05 0.590000 5.473327e-05 0.600000 5.492829e-05 
+ 0.610000 5.511768e-05 0.620000 5.530114e-05 0.630000 5.547797e-05 
+ 0.640000 5.564792e-05 0.650000 5.581025e-05 0.660000 5.596471e-05 
+ 0.670000 5.611085e-05 0.680000 5.624836e-05 0.690000 5.637682e-05 
+ 0.700000 5.649623e-05 0.710000 5.660623e-05 0.720000 5.670677e-05 
+ 0.730000 5.679771e-05 0.740000 5.687916e-05 0.750000 5.695124e-05 
+ 0.760000 5.701383e-05 0.770000 5.706714e-05 0.780000 5.711147e-05 
+ 0.790000 5.714699e-05 0.800000 5.717369e-05)
r_load_0p6900 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.7400) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.7400V
.param vg_value = 0.7400
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.740000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p7400 0 d pwl(0.010000 2.335485e-06 0.020000 4.632619e-06 0.030000 6.889738e-06 
+ 0.040000 9.105194e-06 0.050000 1.127743e-05 0.060000 1.340487e-05 
+ 0.070000 1.548603e-05 0.080000 1.751944e-05 0.090000 1.950375e-05 
+ 0.100000 2.143771e-05 0.110000 2.332002e-05 0.120000 2.514956e-05 
+ 0.130000 2.692530e-05 0.140000 2.864633e-05 0.150000 3.031175e-05 
+ 0.160000 3.192089e-05 0.170000 3.347315e-05 0.180000 3.496806e-05 
+ 0.190000 3.640526e-05 0.200000 3.778467e-05 0.210000 3.910619e-05 
+ 0.220000 4.036998e-05 0.230000 4.157642e-05 0.240000 4.272586e-05 
+ 0.250000 4.381899e-05 0.260000 4.485675e-05 0.270000 4.584006e-05 
+ 0.280000 4.677005e-05 0.290000 4.764822e-05 0.300000 4.847587e-05 
+ 0.310000 4.925497e-05 0.320000 4.998712e-05 0.330000 5.067448e-05 
+ 0.340000 5.131908e-05 0.350000 5.192315e-05 0.360000 5.248910e-05 
+ 0.370000 5.301921e-05 0.380000 5.351596e-05 0.390000 5.398197e-05 
+ 0.400000 5.441961e-05 0.410000 5.483147e-05 0.420000 5.521990e-05 
+ 0.430000 5.558736e-05 0.440000 5.593622e-05 0.450000 5.626845e-05 
+ 0.460000 5.658625e-05 0.470000 5.689164e-05 0.480000 5.718620e-05 
+ 0.490000 5.747164e-05 0.500000 5.774921e-05 0.510000 5.802029e-05 
+ 0.520000 5.828557e-05 0.530000 5.854610e-05 0.540000 5.880238e-05 
+ 0.550000 5.905479e-05 0.560000 5.930361e-05 0.570000 5.954886e-05 
+ 0.580000 5.979034e-05 0.590000 6.002801e-05 0.600000 6.026149e-05 
+ 0.610000 6.049020e-05 0.620000 6.071377e-05 0.630000 6.093162e-05 
+ 0.640000 6.114311e-05 0.650000 6.134756e-05 0.660000 6.154446e-05 
+ 0.670000 6.173318e-05 0.680000 6.191316e-05 0.690000 6.208404e-05 
+ 0.700000 6.224509e-05 0.710000 6.239603e-05 0.720000 6.253648e-05 
+ 0.730000 6.266623e-05 0.740000 6.278519e-05 0.750000 6.289294e-05 
+ 0.760000 6.298974e-05 0.770000 6.307541e-05 0.780000 6.315006e-05 
+ 0.790000 6.321379e-05 0.800000 6.326686e-05)
r_load_0p7400 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* DC Sweep - Gate Voltage (Vg=0.8000) and Drain Voltage (Vd)
******************************************************************
* For Vg = 0.8000V
.param vg_value = 0.8000
* Fix gate voltage for this sweep
e_vg_fix g_orig 0 dc = 0.800000
* Create PWL current source based on data from NN model for this Vg
* The format is: Vd1 Id1 Vd2 Id2 Vd3 Id3 etc.
i_pred_0p8000 0 d pwl(0.010000 2.375805e-06 0.020000 4.716832e-06 0.030000 7.021654e-06 
+ 0.040000 9.288861e-06 0.050000 1.151707e-05 0.060000 1.370497e-05 
+ 0.070000 1.585118e-05 0.080000 1.795450e-05 0.090000 2.001362e-05 
+ 0.100000 2.202743e-05 0.110000 2.399474e-05 0.120000 2.591446e-05 
+ 0.130000 2.778564e-05 0.140000 2.960726e-05 0.150000 3.137843e-05 
+ 0.160000 3.309840e-05 0.170000 3.476649e-05 0.180000 3.638191e-05 
+ 0.190000 3.794425e-05 0.200000 3.945306e-05 0.210000 4.090800e-05 
+ 0.220000 4.230891e-05 0.230000 4.365565e-05 0.240000 4.494823e-05 
+ 0.250000 4.618688e-05 0.260000 4.737185e-05 0.270000 4.850364e-05 
+ 0.280000 4.958295e-05 0.290000 5.061038e-05 0.300000 5.158685e-05 
+ 0.310000 5.251346e-05 0.320000 5.339147e-05 0.330000 5.422210e-05 
+ 0.340000 5.500690e-05 0.350000 5.574755e-05 0.360000 5.644592e-05 
+ 0.370000 5.710366e-05 0.380000 5.772306e-05 0.390000 5.830600e-05 
+ 0.400000 5.885476e-05 0.410000 5.937148e-05 0.420000 5.985878e-05 
+ 0.430000 6.031862e-05 0.440000 6.075341e-05 0.450000 6.116562e-05 
+ 0.460000 6.155744e-05 0.470000 6.193099e-05 0.480000 6.228840e-05 
+ 0.490000 6.263168e-05 0.500000 6.296250e-05 0.510000 6.328297e-05 
+ 0.520000 6.359438e-05 0.530000 6.389826e-05 0.540000 6.419554e-05 
+ 0.550000 6.448752e-05 0.560000 6.477468e-05 0.570000 6.505780e-05 
+ 0.580000 6.533727e-05 0.590000 6.561325e-05 0.600000 6.588591e-05 
+ 0.610000 6.615490e-05 0.620000 6.642012e-05 0.630000 6.668107e-05 
+ 0.640000 6.693742e-05 0.650000 6.718834e-05 0.660000 6.743318e-05 
+ 0.670000 6.767150e-05 0.680000 6.790227e-05 0.690000 6.812488e-05 
+ 0.700000 6.833874e-05 0.710000 6.854282e-05 0.720000 6.873689e-05 
+ 0.730000 6.892017e-05 0.740000 6.909197e-05 0.750000 6.925234e-05 
+ 0.760000 6.940035e-05 0.770000 6.953610e-05 0.780000 6.965944e-05 
+ 0.790000 6.976999e-05 0.800000 6.986799e-05)
r_load_0p8000 d 0 1e6
* Run DC sweep
.dc vd 0 0.8 0.01

******************************************************************
* Probe Statements
******************************************************************
* Probe the gate voltage
.probe dc v(g_orig)

* Probe the drain voltage
.probe dc v(d)

* Probe the actual MOSFET drain current
.probe dc i(vd_orig)

* Probe the predicted (neural network) currents
.probe dc i(i_pred_0p0100)
.probe dc i(i_pred_0p0600)
.probe dc i(i_pred_0p1100)
.probe dc i(i_pred_0p1600)
.probe dc i(i_pred_0p2200)
.probe dc i(i_pred_0p2700)
.probe dc i(i_pred_0p3200)
.probe dc i(i_pred_0p3700)
.probe dc i(i_pred_0p4300)
.probe dc i(i_pred_0p4800)
.probe dc i(i_pred_0p5300)
.probe dc i(i_pred_0p5800)
.probe dc i(i_pred_0p6400)
.probe dc i(i_pred_0p6900)
.probe dc i(i_pred_0p7400)
.probe dc i(i_pred_0p8000)

* Additional options
.option post=2 measout

.end
